library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom2 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"7c3c0000",
     1 => x"7c7c4040",
     2 => x"3c1c0000",
     3 => x"1c3c6060",
     4 => x"607c3c00",
     5 => x"3c7c6030",
     6 => x"386c4400",
     7 => x"446c3810",
     8 => x"bc1c0000",
     9 => x"1c3c60e0",
    10 => x"64440000",
    11 => x"444c5c74",
    12 => x"08080000",
    13 => x"4141773e",
    14 => x"00000000",
    15 => x"00007f7f",
    16 => x"41410000",
    17 => x"08083e77",
    18 => x"01010200",
    19 => x"01020203",
    20 => x"7f7f7f00",
    21 => x"7f7f7f7f",
    22 => x"1c080800",
    23 => x"7f3e3e1c",
    24 => x"3e7f7f7f",
    25 => x"081c1c3e",
    26 => x"18100008",
    27 => x"10187c7c",
    28 => x"30100000",
    29 => x"10307c7c",
    30 => x"60301000",
    31 => x"061e7860",
    32 => x"3c664200",
    33 => x"42663c18",
    34 => x"6a387800",
    35 => x"386cc6c2",
    36 => x"00006000",
    37 => x"60000060",
    38 => x"5b5e0e00",
    39 => x"1e0e5d5c",
    40 => x"ecc24c71",
    41 => x"c04dbfd5",
    42 => x"741ec04b",
    43 => x"87c702ab",
    44 => x"c048a6c4",
    45 => x"c487c578",
    46 => x"78c148a6",
    47 => x"731e66c4",
    48 => x"87dfee49",
    49 => x"e0c086c8",
    50 => x"87eeef49",
    51 => x"6a4aa5c4",
    52 => x"87f0f049",
    53 => x"cb87c6f1",
    54 => x"c883c185",
    55 => x"ff04abb7",
    56 => x"262687c7",
    57 => x"264c264d",
    58 => x"1e4f264b",
    59 => x"ecc24a71",
    60 => x"ecc25ad9",
    61 => x"78c748d9",
    62 => x"87ddfe49",
    63 => x"731e4f26",
    64 => x"c04a711e",
    65 => x"d303aab7",
    66 => x"f7d2c287",
    67 => x"87c405bf",
    68 => x"87c24bc1",
    69 => x"d2c24bc0",
    70 => x"87c45bfb",
    71 => x"5afbd2c2",
    72 => x"bff7d2c2",
    73 => x"c19ac14a",
    74 => x"ec49a2c0",
    75 => x"48fc87e8",
    76 => x"bff7d2c2",
    77 => x"87effe78",
    78 => x"c44a711e",
    79 => x"49721e66",
    80 => x"2687f9ea",
    81 => x"711e4f26",
    82 => x"48d4ff4a",
    83 => x"ff78ffc3",
    84 => x"e1c048d0",
    85 => x"48d4ff78",
    86 => x"497278c1",
    87 => x"787131c4",
    88 => x"c048d0ff",
    89 => x"4f2678e0",
    90 => x"5c5b5e0e",
    91 => x"86f40e5d",
    92 => x"c048a6c4",
    93 => x"bfec4b78",
    94 => x"d5ecc27e",
    95 => x"bfe84dbf",
    96 => x"f7d2c24c",
    97 => x"fee249bf",
    98 => x"49eecb87",
    99 => x"cc87f0cc",
   100 => x"49c758a6",
   101 => x"7087f3e6",
   102 => x"87c80598",
   103 => x"99c1496e",
   104 => x"87c3c102",
   105 => x"bfec4bc1",
   106 => x"f7d2c27e",
   107 => x"d6e249bf",
   108 => x"4966c887",
   109 => x"7087d4cc",
   110 => x"87d80298",
   111 => x"bfefd2c2",
   112 => x"c2b9c149",
   113 => x"7159f3d2",
   114 => x"cb87fbfd",
   115 => x"eecb49ee",
   116 => x"58a6cc87",
   117 => x"f1e549c7",
   118 => x"05987087",
   119 => x"6e87c5ff",
   120 => x"0599c149",
   121 => x"7387fdfe",
   122 => x"87d0029b",
   123 => x"cdfc49ff",
   124 => x"49dac187",
   125 => x"c487d3e5",
   126 => x"78c148a6",
   127 => x"bff7d2c2",
   128 => x"87e9c005",
   129 => x"e549fdc3",
   130 => x"fac387c0",
   131 => x"87fae449",
   132 => x"ffc34974",
   133 => x"c01e7199",
   134 => x"87dcfc49",
   135 => x"b7c84974",
   136 => x"c11e7129",
   137 => x"87d0fc49",
   138 => x"ecc886c8",
   139 => x"c3497487",
   140 => x"b7c899ff",
   141 => x"74b4712c",
   142 => x"87dd029c",
   143 => x"bff3d2c2",
   144 => x"87c7ca49",
   145 => x"c4059870",
   146 => x"d24cc087",
   147 => x"49e0c287",
   148 => x"c287ecc9",
   149 => x"c658f7d2",
   150 => x"f3d2c287",
   151 => x"7478c048",
   152 => x"0599c249",
   153 => x"ebc387cd",
   154 => x"87dee349",
   155 => x"99c24970",
   156 => x"c187cf02",
   157 => x"6e7ea5d8",
   158 => x"c5c002bf",
   159 => x"49fb4b87",
   160 => x"49740f73",
   161 => x"cd0599c1",
   162 => x"49f4c387",
   163 => x"7087fbe2",
   164 => x"0299c249",
   165 => x"d8c187cf",
   166 => x"bf6e7ea5",
   167 => x"87c5c002",
   168 => x"7349fa4b",
   169 => x"c849740f",
   170 => x"87ce0599",
   171 => x"e249f5c3",
   172 => x"497087d8",
   173 => x"c00299c2",
   174 => x"ecc287e5",
   175 => x"c002bfd9",
   176 => x"c14887ca",
   177 => x"ddecc288",
   178 => x"87cec058",
   179 => x"4aa5d8c1",
   180 => x"c5c0026a",
   181 => x"49ff4b87",
   182 => x"a6c40f73",
   183 => x"7478c148",
   184 => x"0599c449",
   185 => x"c387cec0",
   186 => x"dde149f2",
   187 => x"c2497087",
   188 => x"ecc00299",
   189 => x"d9ecc287",
   190 => x"c7487ebf",
   191 => x"c003a8b7",
   192 => x"486e87cb",
   193 => x"ecc280c1",
   194 => x"cfc058dd",
   195 => x"a5d8c187",
   196 => x"02bf6e7e",
   197 => x"4b87c5c0",
   198 => x"0f7349fe",
   199 => x"c148a6c4",
   200 => x"49fdc378",
   201 => x"7087e3e0",
   202 => x"0299c249",
   203 => x"c287e5c0",
   204 => x"02bfd9ec",
   205 => x"c287c9c0",
   206 => x"c048d9ec",
   207 => x"87cfc078",
   208 => x"7ea5d8c1",
   209 => x"c002bf6e",
   210 => x"fd4b87c5",
   211 => x"c40f7349",
   212 => x"78c148a6",
   213 => x"ff49fac3",
   214 => x"7087efdf",
   215 => x"0299c249",
   216 => x"c287e9c0",
   217 => x"48bfd9ec",
   218 => x"03a8b7c7",
   219 => x"c287c9c0",
   220 => x"c748d9ec",
   221 => x"87cfc078",
   222 => x"7ea5d8c1",
   223 => x"c002bf6e",
   224 => x"fc4b87c5",
   225 => x"c40f7349",
   226 => x"78c148a6",
   227 => x"ecc24bc0",
   228 => x"50c048d4",
   229 => x"c449eecb",
   230 => x"a6cc87e5",
   231 => x"d4ecc258",
   232 => x"c105bf97",
   233 => x"497487de",
   234 => x"0599f0c3",
   235 => x"c187cdc0",
   236 => x"deff49da",
   237 => x"987087d4",
   238 => x"87c8c102",
   239 => x"bfe84bc1",
   240 => x"ffc3494c",
   241 => x"2cb7c899",
   242 => x"d2c2b471",
   243 => x"ff49bff7",
   244 => x"c887f4d9",
   245 => x"f2c34966",
   246 => x"02987087",
   247 => x"c287c6c0",
   248 => x"c148d4ec",
   249 => x"d4ecc250",
   250 => x"c005bf97",
   251 => x"497487d6",
   252 => x"0599f0c3",
   253 => x"c187c5ff",
   254 => x"ddff49da",
   255 => x"987087cc",
   256 => x"87f8fe05",
   257 => x"c0029b73",
   258 => x"a6c887dc",
   259 => x"d9ecc248",
   260 => x"66c878bf",
   261 => x"7591cb49",
   262 => x"bf6e7ea1",
   263 => x"87c6c002",
   264 => x"4966c84b",
   265 => x"66c40f73",
   266 => x"87c8c002",
   267 => x"bfd9ecc2",
   268 => x"87e5f149",
   269 => x"bffbd2c2",
   270 => x"87ddc002",
   271 => x"87cbc249",
   272 => x"c0029870",
   273 => x"ecc287d3",
   274 => x"f149bfd9",
   275 => x"49c087cb",
   276 => x"c287ebf2",
   277 => x"c048fbd2",
   278 => x"f28ef478",
   279 => x"5e0e87c5",
   280 => x"0e5d5c5b",
   281 => x"c24c711e",
   282 => x"49bfd5ec",
   283 => x"4da1cdc1",
   284 => x"6981d1c1",
   285 => x"029c747e",
   286 => x"a5c487cf",
   287 => x"c27b744b",
   288 => x"49bfd5ec",
   289 => x"6e87e4f1",
   290 => x"059c747b",
   291 => x"4bc087c4",
   292 => x"4bc187c2",
   293 => x"e5f14973",
   294 => x"0266d487",
   295 => x"de4987c7",
   296 => x"c24a7087",
   297 => x"c24ac087",
   298 => x"265affd2",
   299 => x"0087f4f0",
   300 => x"00000000",
   301 => x"00000000",
   302 => x"00000000",
   303 => x"1e000000",
   304 => x"c8ff4a71",
   305 => x"a17249bf",
   306 => x"1e4f2648",
   307 => x"89bfc8ff",
   308 => x"c0c0c0fe",
   309 => x"01a9c0c0",
   310 => x"4ac087c4",
   311 => x"4ac187c2",
   312 => x"4f264872",
   313 => x"5c5b5e0e",
   314 => x"4b710e5d",
   315 => x"d04cd4ff",
   316 => x"78c04866",
   317 => x"dbff49d6",
   318 => x"ffc387c8",
   319 => x"c3496c7c",
   320 => x"4d7199ff",
   321 => x"99f0c349",
   322 => x"05a9e0c1",
   323 => x"ffc387cb",
   324 => x"c3486c7c",
   325 => x"0866d098",
   326 => x"7cffc378",
   327 => x"c8494a6c",
   328 => x"7cffc331",
   329 => x"b2714a6c",
   330 => x"31c84972",
   331 => x"6c7cffc3",
   332 => x"72b2714a",
   333 => x"c331c849",
   334 => x"4a6c7cff",
   335 => x"d0ffb271",
   336 => x"78e0c048",
   337 => x"c2029b73",
   338 => x"757b7287",
   339 => x"264d2648",
   340 => x"264b264c",
   341 => x"4f261e4f",
   342 => x"5c5b5e0e",
   343 => x"7686f80e",
   344 => x"49a6c81e",
   345 => x"c487fdfd",
   346 => x"6e4b7086",
   347 => x"03a8c248",
   348 => x"7387f0c2",
   349 => x"9af0c34a",
   350 => x"02aad0c1",
   351 => x"e0c187c7",
   352 => x"dec205aa",
   353 => x"c8497387",
   354 => x"87c30299",
   355 => x"7387c6ff",
   356 => x"c29cc34c",
   357 => x"c2c105ac",
   358 => x"4966c487",
   359 => x"1e7131c9",
   360 => x"d44a66c4",
   361 => x"ddecc292",
   362 => x"fe817249",
   363 => x"d887d4d0",
   364 => x"cdd8ff49",
   365 => x"1ec0c887",
   366 => x"49c6dbc2",
   367 => x"87deecfd",
   368 => x"c048d0ff",
   369 => x"dbc278e0",
   370 => x"66cc1ec6",
   371 => x"c292d44a",
   372 => x"7249ddec",
   373 => x"dccefe81",
   374 => x"c186cc87",
   375 => x"c2c105ac",
   376 => x"4966c487",
   377 => x"1e7131c9",
   378 => x"d44a66c4",
   379 => x"ddecc292",
   380 => x"fe817249",
   381 => x"c287cccf",
   382 => x"c81ec6db",
   383 => x"92d44a66",
   384 => x"49ddecc2",
   385 => x"ccfe8172",
   386 => x"49d787dd",
   387 => x"87f2d6ff",
   388 => x"c21ec0c8",
   389 => x"fd49c6db",
   390 => x"cc87dcea",
   391 => x"48d0ff86",
   392 => x"f878e0c0",
   393 => x"87e7fc8e",
   394 => x"5c5b5e0e",
   395 => x"4a710e5d",
   396 => x"d04cd4ff",
   397 => x"b7c34d66",
   398 => x"87c506ad",
   399 => x"dac148c0",
   400 => x"751e7287",
   401 => x"c293d44b",
   402 => x"7383ddec",
   403 => x"e4c6fe49",
   404 => x"6b83c887",
   405 => x"48d0ff4b",
   406 => x"dd78e1c8",
   407 => x"c349737c",
   408 => x"7c7199ff",
   409 => x"b7c84973",
   410 => x"99ffc329",
   411 => x"49737c71",
   412 => x"c329b7d0",
   413 => x"7c7199ff",
   414 => x"b7d84973",
   415 => x"c07c7129",
   416 => x"7c7c7c7c",
   417 => x"7c7c7c7c",
   418 => x"7c7c7c7c",
   419 => x"7578e0c0",
   420 => x"ff49dc1e",
   421 => x"c887d0d5",
   422 => x"fa487386",
   423 => x"fa4887ef",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
