
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom1 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom1 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"c8",x"ed",x"c2",x"87"),
    12 => (x"86",x"c0",x"c8",x"4e"),
    13 => (x"49",x"c8",x"ed",x"c2"),
    14 => (x"48",x"e0",x"da",x"c2"),
    15 => (x"40",x"40",x"c0",x"89"),
    16 => (x"89",x"d0",x"40",x"40"),
    17 => (x"c1",x"87",x"f6",x"03"),
    18 => (x"00",x"87",x"c3",x"e2"),
    19 => (x"72",x"1e",x"87",x"fd"),
    20 => (x"12",x"1e",x"73",x"1e"),
    21 => (x"ca",x"02",x"11",x"48"),
    22 => (x"df",x"c3",x"4b",x"87"),
    23 => (x"88",x"73",x"9b",x"98"),
    24 => (x"26",x"87",x"f0",x"02"),
    25 => (x"26",x"4a",x"26",x"4b"),
    26 => (x"1e",x"73",x"1e",x"4f"),
    27 => (x"8b",x"c1",x"1e",x"72"),
    28 => (x"12",x"87",x"ca",x"04"),
    29 => (x"c4",x"02",x"11",x"48"),
    30 => (x"f1",x"02",x"88",x"87"),
    31 => (x"26",x"4a",x"26",x"87"),
    32 => (x"1e",x"4f",x"26",x"4b"),
    33 => (x"1e",x"73",x"1e",x"74"),
    34 => (x"8b",x"c1",x"1e",x"72"),
    35 => (x"12",x"87",x"d0",x"04"),
    36 => (x"ca",x"02",x"11",x"48"),
    37 => (x"df",x"c3",x"4c",x"87"),
    38 => (x"88",x"74",x"9c",x"98"),
    39 => (x"26",x"87",x"eb",x"02"),
    40 => (x"26",x"4b",x"26",x"4a"),
    41 => (x"1e",x"4f",x"26",x"4c"),
    42 => (x"73",x"81",x"48",x"73"),
    43 => (x"87",x"c5",x"02",x"a9"),
    44 => (x"f6",x"05",x"53",x"12"),
    45 => (x"1e",x"4f",x"26",x"87"),
    46 => (x"66",x"c4",x"4a",x"71"),
    47 => (x"88",x"c1",x"48",x"49"),
    48 => (x"71",x"58",x"a6",x"c8"),
    49 => (x"87",x"d4",x"02",x"99"),
    50 => (x"d4",x"ff",x"48",x"12"),
    51 => (x"66",x"c4",x"78",x"08"),
    52 => (x"88",x"c1",x"48",x"49"),
    53 => (x"71",x"58",x"a6",x"c8"),
    54 => (x"87",x"ec",x"05",x"99"),
    55 => (x"71",x"1e",x"4f",x"26"),
    56 => (x"49",x"66",x"c4",x"4a"),
    57 => (x"c8",x"88",x"c1",x"48"),
    58 => (x"99",x"71",x"58",x"a6"),
    59 => (x"ff",x"87",x"d6",x"02"),
    60 => (x"ff",x"c3",x"48",x"d4"),
    61 => (x"c4",x"52",x"68",x"78"),
    62 => (x"c1",x"48",x"49",x"66"),
    63 => (x"58",x"a6",x"c8",x"88"),
    64 => (x"ea",x"05",x"99",x"71"),
    65 => (x"1e",x"4f",x"26",x"87"),
    66 => (x"d4",x"ff",x"1e",x"73"),
    67 => (x"7b",x"ff",x"c3",x"4b"),
    68 => (x"ff",x"c3",x"4a",x"6b"),
    69 => (x"c8",x"49",x"6b",x"7b"),
    70 => (x"c3",x"b1",x"72",x"32"),
    71 => (x"4a",x"6b",x"7b",x"ff"),
    72 => (x"b2",x"71",x"31",x"c8"),
    73 => (x"6b",x"7b",x"ff",x"c3"),
    74 => (x"72",x"32",x"c8",x"49"),
    75 => (x"c4",x"48",x"71",x"b1"),
    76 => (x"26",x"4d",x"26",x"87"),
    77 => (x"26",x"4b",x"26",x"4c"),
    78 => (x"5b",x"5e",x"0e",x"4f"),
    79 => (x"71",x"0e",x"5d",x"5c"),
    80 => (x"4c",x"d4",x"ff",x"4a"),
    81 => (x"ff",x"c3",x"48",x"72"),
    82 => (x"c2",x"7c",x"70",x"98"),
    83 => (x"05",x"bf",x"e0",x"da"),
    84 => (x"66",x"d0",x"87",x"c8"),
    85 => (x"d4",x"30",x"c9",x"48"),
    86 => (x"66",x"d0",x"58",x"a6"),
    87 => (x"71",x"29",x"d8",x"49"),
    88 => (x"98",x"ff",x"c3",x"48"),
    89 => (x"66",x"d0",x"7c",x"70"),
    90 => (x"c3",x"29",x"d0",x"49"),
    91 => (x"7c",x"71",x"99",x"ff"),
    92 => (x"c8",x"49",x"66",x"d0"),
    93 => (x"99",x"ff",x"c3",x"29"),
    94 => (x"66",x"d0",x"7c",x"71"),
    95 => (x"99",x"ff",x"c3",x"49"),
    96 => (x"49",x"72",x"7c",x"71"),
    97 => (x"48",x"71",x"29",x"d0"),
    98 => (x"70",x"98",x"ff",x"c3"),
    99 => (x"c9",x"4b",x"6c",x"7c"),
   100 => (x"c3",x"4d",x"ff",x"f0"),
   101 => (x"d0",x"05",x"ab",x"ff"),
   102 => (x"7c",x"ff",x"c3",x"87"),
   103 => (x"8d",x"c1",x"4b",x"6c"),
   104 => (x"c3",x"87",x"c6",x"02"),
   105 => (x"f0",x"02",x"ab",x"ff"),
   106 => (x"fe",x"48",x"73",x"87"),
   107 => (x"c0",x"1e",x"87",x"c3"),
   108 => (x"48",x"d4",x"ff",x"49"),
   109 => (x"c1",x"78",x"ff",x"c3"),
   110 => (x"b7",x"c8",x"c3",x"81"),
   111 => (x"87",x"f1",x"04",x"a9"),
   112 => (x"73",x"1e",x"4f",x"26"),
   113 => (x"c4",x"87",x"e7",x"1e"),
   114 => (x"c0",x"4b",x"df",x"f8"),
   115 => (x"f0",x"ff",x"c0",x"1e"),
   116 => (x"fd",x"49",x"f7",x"c1"),
   117 => (x"86",x"c4",x"87",x"e3"),
   118 => (x"c0",x"05",x"a8",x"c1"),
   119 => (x"d4",x"ff",x"87",x"ea"),
   120 => (x"78",x"ff",x"c3",x"48"),
   121 => (x"c0",x"c0",x"c0",x"c1"),
   122 => (x"c0",x"1e",x"c0",x"c0"),
   123 => (x"e9",x"c1",x"f0",x"e1"),
   124 => (x"87",x"c5",x"fd",x"49"),
   125 => (x"98",x"70",x"86",x"c4"),
   126 => (x"ff",x"87",x"ca",x"05"),
   127 => (x"ff",x"c3",x"48",x"d4"),
   128 => (x"cb",x"48",x"c1",x"78"),
   129 => (x"87",x"e6",x"fe",x"87"),
   130 => (x"fe",x"05",x"8b",x"c1"),
   131 => (x"48",x"c0",x"87",x"fd"),
   132 => (x"1e",x"87",x"e2",x"fc"),
   133 => (x"d4",x"ff",x"1e",x"73"),
   134 => (x"78",x"ff",x"c3",x"48"),
   135 => (x"1e",x"c0",x"4b",x"d3"),
   136 => (x"c1",x"f0",x"ff",x"c0"),
   137 => (x"d0",x"fc",x"49",x"c1"),
   138 => (x"70",x"86",x"c4",x"87"),
   139 => (x"87",x"ca",x"05",x"98"),
   140 => (x"c3",x"48",x"d4",x"ff"),
   141 => (x"48",x"c1",x"78",x"ff"),
   142 => (x"f1",x"fd",x"87",x"cb"),
   143 => (x"05",x"8b",x"c1",x"87"),
   144 => (x"c0",x"87",x"db",x"ff"),
   145 => (x"87",x"ed",x"fb",x"48"),
   146 => (x"5c",x"5b",x"5e",x"0e"),
   147 => (x"4c",x"d4",x"ff",x"0e"),
   148 => (x"c6",x"87",x"db",x"fd"),
   149 => (x"e1",x"c0",x"1e",x"ea"),
   150 => (x"49",x"c8",x"c1",x"f0"),
   151 => (x"c4",x"87",x"da",x"fb"),
   152 => (x"02",x"a8",x"c1",x"86"),
   153 => (x"ea",x"fe",x"87",x"c8"),
   154 => (x"c1",x"48",x"c0",x"87"),
   155 => (x"d6",x"fa",x"87",x"e2"),
   156 => (x"cf",x"49",x"70",x"87"),
   157 => (x"c6",x"99",x"ff",x"ff"),
   158 => (x"c8",x"02",x"a9",x"ea"),
   159 => (x"87",x"d3",x"fe",x"87"),
   160 => (x"cb",x"c1",x"48",x"c0"),
   161 => (x"7c",x"ff",x"c3",x"87"),
   162 => (x"fc",x"4b",x"f1",x"c0"),
   163 => (x"98",x"70",x"87",x"f4"),
   164 => (x"87",x"eb",x"c0",x"02"),
   165 => (x"ff",x"c0",x"1e",x"c0"),
   166 => (x"49",x"fa",x"c1",x"f0"),
   167 => (x"c4",x"87",x"da",x"fa"),
   168 => (x"05",x"98",x"70",x"86"),
   169 => (x"ff",x"c3",x"87",x"d9"),
   170 => (x"c3",x"49",x"6c",x"7c"),
   171 => (x"7c",x"7c",x"7c",x"ff"),
   172 => (x"99",x"c0",x"c1",x"7c"),
   173 => (x"c1",x"87",x"c4",x"02"),
   174 => (x"c0",x"87",x"d5",x"48"),
   175 => (x"c2",x"87",x"d1",x"48"),
   176 => (x"87",x"c4",x"05",x"ab"),
   177 => (x"87",x"c8",x"48",x"c0"),
   178 => (x"fe",x"05",x"8b",x"c1"),
   179 => (x"48",x"c0",x"87",x"fd"),
   180 => (x"1e",x"87",x"e0",x"f9"),
   181 => (x"da",x"c2",x"1e",x"73"),
   182 => (x"78",x"c1",x"48",x"e0"),
   183 => (x"d0",x"ff",x"4b",x"c7"),
   184 => (x"fb",x"78",x"c2",x"48"),
   185 => (x"d0",x"ff",x"87",x"c8"),
   186 => (x"c0",x"78",x"c3",x"48"),
   187 => (x"d0",x"e5",x"c0",x"1e"),
   188 => (x"f9",x"49",x"c0",x"c1"),
   189 => (x"86",x"c4",x"87",x"c3"),
   190 => (x"c1",x"05",x"a8",x"c1"),
   191 => (x"ab",x"c2",x"4b",x"87"),
   192 => (x"c0",x"87",x"c5",x"05"),
   193 => (x"87",x"f9",x"c0",x"48"),
   194 => (x"ff",x"05",x"8b",x"c1"),
   195 => (x"f7",x"fc",x"87",x"d0"),
   196 => (x"e4",x"da",x"c2",x"87"),
   197 => (x"05",x"98",x"70",x"58"),
   198 => (x"1e",x"c1",x"87",x"cd"),
   199 => (x"c1",x"f0",x"ff",x"c0"),
   200 => (x"d4",x"f8",x"49",x"d0"),
   201 => (x"ff",x"86",x"c4",x"87"),
   202 => (x"ff",x"c3",x"48",x"d4"),
   203 => (x"87",x"dd",x"c4",x"78"),
   204 => (x"58",x"e8",x"da",x"c2"),
   205 => (x"c2",x"48",x"d0",x"ff"),
   206 => (x"48",x"d4",x"ff",x"78"),
   207 => (x"c1",x"78",x"ff",x"c3"),
   208 => (x"87",x"f1",x"f7",x"48"),
   209 => (x"5c",x"5b",x"5e",x"0e"),
   210 => (x"4a",x"71",x"0e",x"5d"),
   211 => (x"ff",x"4d",x"ff",x"c3"),
   212 => (x"7c",x"75",x"4c",x"d4"),
   213 => (x"c4",x"48",x"d0",x"ff"),
   214 => (x"7c",x"75",x"78",x"c3"),
   215 => (x"ff",x"c0",x"1e",x"72"),
   216 => (x"49",x"d8",x"c1",x"f0"),
   217 => (x"c4",x"87",x"d2",x"f7"),
   218 => (x"02",x"98",x"70",x"86"),
   219 => (x"48",x"c1",x"87",x"c5"),
   220 => (x"75",x"87",x"ee",x"c0"),
   221 => (x"7c",x"fe",x"c3",x"7c"),
   222 => (x"d4",x"1e",x"c0",x"c8"),
   223 => (x"f6",x"f4",x"49",x"66"),
   224 => (x"75",x"86",x"c4",x"87"),
   225 => (x"75",x"7c",x"75",x"7c"),
   226 => (x"e0",x"da",x"d8",x"7c"),
   227 => (x"6c",x"7c",x"75",x"4b"),
   228 => (x"c1",x"87",x"c5",x"05"),
   229 => (x"87",x"f5",x"05",x"8b"),
   230 => (x"d0",x"ff",x"7c",x"75"),
   231 => (x"c0",x"78",x"c2",x"48"),
   232 => (x"87",x"cd",x"f6",x"48"),
   233 => (x"5c",x"5b",x"5e",x"0e"),
   234 => (x"4b",x"71",x"0e",x"5d"),
   235 => (x"ee",x"c5",x"4c",x"c0"),
   236 => (x"ff",x"4a",x"df",x"cd"),
   237 => (x"ff",x"c3",x"48",x"d4"),
   238 => (x"c3",x"48",x"68",x"78"),
   239 => (x"c0",x"05",x"a8",x"fe"),
   240 => (x"d4",x"ff",x"87",x"fe"),
   241 => (x"02",x"9b",x"73",x"4d"),
   242 => (x"66",x"d0",x"87",x"cc"),
   243 => (x"f4",x"49",x"73",x"1e"),
   244 => (x"86",x"c4",x"87",x"cc"),
   245 => (x"d0",x"ff",x"87",x"d6"),
   246 => (x"78",x"d1",x"c4",x"48"),
   247 => (x"d0",x"7d",x"ff",x"c3"),
   248 => (x"88",x"c1",x"48",x"66"),
   249 => (x"70",x"58",x"a6",x"d4"),
   250 => (x"87",x"f0",x"05",x"98"),
   251 => (x"c3",x"48",x"d4",x"ff"),
   252 => (x"73",x"78",x"78",x"ff"),
   253 => (x"87",x"c5",x"05",x"9b"),
   254 => (x"d0",x"48",x"d0",x"ff"),
   255 => (x"4c",x"4a",x"c1",x"78"),
   256 => (x"fe",x"05",x"8a",x"c1"),
   257 => (x"48",x"74",x"87",x"ed"),
   258 => (x"1e",x"87",x"e6",x"f4"),
   259 => (x"4a",x"71",x"1e",x"73"),
   260 => (x"d4",x"ff",x"4b",x"c0"),
   261 => (x"78",x"ff",x"c3",x"48"),
   262 => (x"c4",x"48",x"d0",x"ff"),
   263 => (x"d4",x"ff",x"78",x"c3"),
   264 => (x"78",x"ff",x"c3",x"48"),
   265 => (x"ff",x"c0",x"1e",x"72"),
   266 => (x"49",x"d1",x"c1",x"f0"),
   267 => (x"c4",x"87",x"ca",x"f4"),
   268 => (x"05",x"98",x"70",x"86"),
   269 => (x"c0",x"c8",x"87",x"d2"),
   270 => (x"49",x"66",x"cc",x"1e"),
   271 => (x"c4",x"87",x"e5",x"fd"),
   272 => (x"ff",x"4b",x"70",x"86"),
   273 => (x"78",x"c2",x"48",x"d0"),
   274 => (x"e8",x"f3",x"48",x"73"),
   275 => (x"5b",x"5e",x"0e",x"87"),
   276 => (x"c0",x"0e",x"5d",x"5c"),
   277 => (x"f0",x"ff",x"c0",x"1e"),
   278 => (x"f3",x"49",x"c9",x"c1"),
   279 => (x"1e",x"d2",x"87",x"db"),
   280 => (x"49",x"e8",x"da",x"c2"),
   281 => (x"c8",x"87",x"fd",x"fc"),
   282 => (x"c1",x"4c",x"c0",x"86"),
   283 => (x"ac",x"b7",x"d2",x"84"),
   284 => (x"c2",x"87",x"f8",x"04"),
   285 => (x"bf",x"97",x"e8",x"da"),
   286 => (x"99",x"c0",x"c3",x"49"),
   287 => (x"05",x"a9",x"c0",x"c1"),
   288 => (x"c2",x"87",x"e7",x"c0"),
   289 => (x"bf",x"97",x"ef",x"da"),
   290 => (x"c2",x"31",x"d0",x"49"),
   291 => (x"bf",x"97",x"f0",x"da"),
   292 => (x"72",x"32",x"c8",x"4a"),
   293 => (x"f1",x"da",x"c2",x"b1"),
   294 => (x"b1",x"4a",x"bf",x"97"),
   295 => (x"ff",x"cf",x"4c",x"71"),
   296 => (x"c1",x"9c",x"ff",x"ff"),
   297 => (x"c1",x"34",x"ca",x"84"),
   298 => (x"da",x"c2",x"87",x"e7"),
   299 => (x"49",x"bf",x"97",x"f1"),
   300 => (x"99",x"c6",x"31",x"c1"),
   301 => (x"97",x"f2",x"da",x"c2"),
   302 => (x"b7",x"c7",x"4a",x"bf"),
   303 => (x"c2",x"b1",x"72",x"2a"),
   304 => (x"bf",x"97",x"ed",x"da"),
   305 => (x"9d",x"cf",x"4d",x"4a"),
   306 => (x"97",x"ee",x"da",x"c2"),
   307 => (x"9a",x"c3",x"4a",x"bf"),
   308 => (x"da",x"c2",x"32",x"ca"),
   309 => (x"4b",x"bf",x"97",x"ef"),
   310 => (x"b2",x"73",x"33",x"c2"),
   311 => (x"97",x"f0",x"da",x"c2"),
   312 => (x"c0",x"c3",x"4b",x"bf"),
   313 => (x"2b",x"b7",x"c6",x"9b"),
   314 => (x"81",x"c2",x"b2",x"73"),
   315 => (x"30",x"71",x"48",x"c1"),
   316 => (x"48",x"c1",x"49",x"70"),
   317 => (x"4d",x"70",x"30",x"75"),
   318 => (x"84",x"c1",x"4c",x"72"),
   319 => (x"c0",x"c8",x"94",x"71"),
   320 => (x"cc",x"06",x"ad",x"b7"),
   321 => (x"b7",x"34",x"c1",x"87"),
   322 => (x"b7",x"c0",x"c8",x"2d"),
   323 => (x"f4",x"ff",x"01",x"ad"),
   324 => (x"f0",x"48",x"74",x"87"),
   325 => (x"5e",x"0e",x"87",x"db"),
   326 => (x"0e",x"5d",x"5c",x"5b"),
   327 => (x"e3",x"c2",x"86",x"f8"),
   328 => (x"78",x"c0",x"48",x"ce"),
   329 => (x"1e",x"c6",x"db",x"c2"),
   330 => (x"de",x"fb",x"49",x"c0"),
   331 => (x"70",x"86",x"c4",x"87"),
   332 => (x"87",x"c5",x"05",x"98"),
   333 => (x"c0",x"c9",x"48",x"c0"),
   334 => (x"c1",x"4d",x"c0",x"87"),
   335 => (x"d9",x"f2",x"c0",x"7e"),
   336 => (x"db",x"c2",x"49",x"bf"),
   337 => (x"c8",x"71",x"4a",x"fc"),
   338 => (x"87",x"dd",x"ec",x"4b"),
   339 => (x"c2",x"05",x"98",x"70"),
   340 => (x"c0",x"7e",x"c0",x"87"),
   341 => (x"49",x"bf",x"d5",x"f2"),
   342 => (x"4a",x"d8",x"dc",x"c2"),
   343 => (x"ec",x"4b",x"c8",x"71"),
   344 => (x"98",x"70",x"87",x"c7"),
   345 => (x"c0",x"87",x"c2",x"05"),
   346 => (x"c0",x"02",x"6e",x"7e"),
   347 => (x"e2",x"c2",x"87",x"fd"),
   348 => (x"c2",x"4d",x"bf",x"cc"),
   349 => (x"bf",x"9f",x"c4",x"e3"),
   350 => (x"d6",x"c5",x"48",x"7e"),
   351 => (x"c7",x"05",x"a8",x"ea"),
   352 => (x"cc",x"e2",x"c2",x"87"),
   353 => (x"87",x"ce",x"4d",x"bf"),
   354 => (x"e9",x"ca",x"48",x"6e"),
   355 => (x"c5",x"02",x"a8",x"d5"),
   356 => (x"c7",x"48",x"c0",x"87"),
   357 => (x"db",x"c2",x"87",x"e3"),
   358 => (x"49",x"75",x"1e",x"c6"),
   359 => (x"c4",x"87",x"ec",x"f9"),
   360 => (x"05",x"98",x"70",x"86"),
   361 => (x"48",x"c0",x"87",x"c5"),
   362 => (x"c0",x"87",x"ce",x"c7"),
   363 => (x"49",x"bf",x"d5",x"f2"),
   364 => (x"4a",x"d8",x"dc",x"c2"),
   365 => (x"ea",x"4b",x"c8",x"71"),
   366 => (x"98",x"70",x"87",x"ef"),
   367 => (x"c2",x"87",x"c8",x"05"),
   368 => (x"c1",x"48",x"ce",x"e3"),
   369 => (x"c0",x"87",x"da",x"78"),
   370 => (x"49",x"bf",x"d9",x"f2"),
   371 => (x"4a",x"fc",x"db",x"c2"),
   372 => (x"ea",x"4b",x"c8",x"71"),
   373 => (x"98",x"70",x"87",x"d3"),
   374 => (x"87",x"c5",x"c0",x"02"),
   375 => (x"d8",x"c6",x"48",x"c0"),
   376 => (x"c4",x"e3",x"c2",x"87"),
   377 => (x"c1",x"49",x"bf",x"97"),
   378 => (x"c0",x"05",x"a9",x"d5"),
   379 => (x"e3",x"c2",x"87",x"cd"),
   380 => (x"49",x"bf",x"97",x"c5"),
   381 => (x"02",x"a9",x"ea",x"c2"),
   382 => (x"c0",x"87",x"c5",x"c0"),
   383 => (x"87",x"f9",x"c5",x"48"),
   384 => (x"97",x"c6",x"db",x"c2"),
   385 => (x"c3",x"48",x"7e",x"bf"),
   386 => (x"c0",x"02",x"a8",x"e9"),
   387 => (x"48",x"6e",x"87",x"ce"),
   388 => (x"02",x"a8",x"eb",x"c3"),
   389 => (x"c0",x"87",x"c5",x"c0"),
   390 => (x"87",x"dd",x"c5",x"48"),
   391 => (x"97",x"d1",x"db",x"c2"),
   392 => (x"05",x"99",x"49",x"bf"),
   393 => (x"c2",x"87",x"cc",x"c0"),
   394 => (x"bf",x"97",x"d2",x"db"),
   395 => (x"02",x"a9",x"c2",x"49"),
   396 => (x"c0",x"87",x"c5",x"c0"),
   397 => (x"87",x"c1",x"c5",x"48"),
   398 => (x"97",x"d3",x"db",x"c2"),
   399 => (x"e3",x"c2",x"48",x"bf"),
   400 => (x"4c",x"70",x"58",x"ca"),
   401 => (x"c2",x"88",x"c1",x"48"),
   402 => (x"c2",x"58",x"ce",x"e3"),
   403 => (x"bf",x"97",x"d4",x"db"),
   404 => (x"c2",x"81",x"75",x"49"),
   405 => (x"bf",x"97",x"d5",x"db"),
   406 => (x"72",x"32",x"c8",x"4a"),
   407 => (x"e7",x"c2",x"7e",x"a1"),
   408 => (x"78",x"6e",x"48",x"db"),
   409 => (x"97",x"d6",x"db",x"c2"),
   410 => (x"a6",x"c8",x"48",x"bf"),
   411 => (x"ce",x"e3",x"c2",x"58"),
   412 => (x"cf",x"c2",x"02",x"bf"),
   413 => (x"d5",x"f2",x"c0",x"87"),
   414 => (x"dc",x"c2",x"49",x"bf"),
   415 => (x"c8",x"71",x"4a",x"d8"),
   416 => (x"87",x"e5",x"e7",x"4b"),
   417 => (x"c0",x"02",x"98",x"70"),
   418 => (x"48",x"c0",x"87",x"c5"),
   419 => (x"c2",x"87",x"ea",x"c3"),
   420 => (x"4c",x"bf",x"c6",x"e3"),
   421 => (x"5c",x"ef",x"e7",x"c2"),
   422 => (x"97",x"eb",x"db",x"c2"),
   423 => (x"31",x"c8",x"49",x"bf"),
   424 => (x"97",x"ea",x"db",x"c2"),
   425 => (x"49",x"a1",x"4a",x"bf"),
   426 => (x"97",x"ec",x"db",x"c2"),
   427 => (x"32",x"d0",x"4a",x"bf"),
   428 => (x"c2",x"49",x"a1",x"72"),
   429 => (x"bf",x"97",x"ed",x"db"),
   430 => (x"72",x"32",x"d8",x"4a"),
   431 => (x"66",x"c4",x"49",x"a1"),
   432 => (x"db",x"e7",x"c2",x"91"),
   433 => (x"e7",x"c2",x"81",x"bf"),
   434 => (x"db",x"c2",x"59",x"e3"),
   435 => (x"4a",x"bf",x"97",x"f3"),
   436 => (x"db",x"c2",x"32",x"c8"),
   437 => (x"4b",x"bf",x"97",x"f2"),
   438 => (x"db",x"c2",x"4a",x"a2"),
   439 => (x"4b",x"bf",x"97",x"f4"),
   440 => (x"a2",x"73",x"33",x"d0"),
   441 => (x"f5",x"db",x"c2",x"4a"),
   442 => (x"cf",x"4b",x"bf",x"97"),
   443 => (x"73",x"33",x"d8",x"9b"),
   444 => (x"e7",x"c2",x"4a",x"a2"),
   445 => (x"8a",x"c2",x"5a",x"e7"),
   446 => (x"e7",x"c2",x"92",x"74"),
   447 => (x"a1",x"72",x"48",x"e7"),
   448 => (x"87",x"c1",x"c1",x"78"),
   449 => (x"97",x"d8",x"db",x"c2"),
   450 => (x"31",x"c8",x"49",x"bf"),
   451 => (x"97",x"d7",x"db",x"c2"),
   452 => (x"49",x"a1",x"4a",x"bf"),
   453 => (x"ff",x"c7",x"31",x"c5"),
   454 => (x"c2",x"29",x"c9",x"81"),
   455 => (x"c2",x"59",x"ef",x"e7"),
   456 => (x"bf",x"97",x"dd",x"db"),
   457 => (x"c2",x"32",x"c8",x"4a"),
   458 => (x"bf",x"97",x"dc",x"db"),
   459 => (x"c4",x"4a",x"a2",x"4b"),
   460 => (x"82",x"6e",x"92",x"66"),
   461 => (x"5a",x"eb",x"e7",x"c2"),
   462 => (x"48",x"e3",x"e7",x"c2"),
   463 => (x"e7",x"c2",x"78",x"c0"),
   464 => (x"a1",x"72",x"48",x"df"),
   465 => (x"ef",x"e7",x"c2",x"78"),
   466 => (x"e3",x"e7",x"c2",x"48"),
   467 => (x"e7",x"c2",x"78",x"bf"),
   468 => (x"e7",x"c2",x"48",x"f3"),
   469 => (x"c2",x"78",x"bf",x"e7"),
   470 => (x"02",x"bf",x"ce",x"e3"),
   471 => (x"74",x"87",x"c9",x"c0"),
   472 => (x"70",x"30",x"c4",x"48"),
   473 => (x"87",x"c9",x"c0",x"7e"),
   474 => (x"bf",x"eb",x"e7",x"c2"),
   475 => (x"70",x"30",x"c4",x"48"),
   476 => (x"d2",x"e3",x"c2",x"7e"),
   477 => (x"c1",x"78",x"6e",x"48"),
   478 => (x"26",x"8e",x"f8",x"48"),
   479 => (x"26",x"4c",x"26",x"4d"),
   480 => (x"0e",x"4f",x"26",x"4b"),
   481 => (x"5d",x"5c",x"5b",x"5e"),
   482 => (x"c2",x"4a",x"71",x"0e"),
   483 => (x"02",x"bf",x"ce",x"e3"),
   484 => (x"4b",x"72",x"87",x"cb"),
   485 => (x"4d",x"72",x"2b",x"c7"),
   486 => (x"c9",x"9d",x"ff",x"c1"),
   487 => (x"c8",x"4b",x"72",x"87"),
   488 => (x"c3",x"4d",x"72",x"2b"),
   489 => (x"e7",x"c2",x"9d",x"ff"),
   490 => (x"c0",x"83",x"bf",x"db"),
   491 => (x"ab",x"bf",x"d1",x"f2"),
   492 => (x"c0",x"87",x"d9",x"02"),
   493 => (x"c2",x"5b",x"d5",x"f2"),
   494 => (x"73",x"1e",x"c6",x"db"),
   495 => (x"87",x"cb",x"f1",x"49"),
   496 => (x"98",x"70",x"86",x"c4"),
   497 => (x"c0",x"87",x"c5",x"05"),
   498 => (x"87",x"e6",x"c0",x"48"),
   499 => (x"bf",x"ce",x"e3",x"c2"),
   500 => (x"75",x"87",x"d2",x"02"),
   501 => (x"c2",x"91",x"c4",x"49"),
   502 => (x"69",x"81",x"c6",x"db"),
   503 => (x"ff",x"ff",x"cf",x"4c"),
   504 => (x"cb",x"9c",x"ff",x"ff"),
   505 => (x"c2",x"49",x"75",x"87"),
   506 => (x"c6",x"db",x"c2",x"91"),
   507 => (x"4c",x"69",x"9f",x"81"),
   508 => (x"c6",x"fe",x"48",x"74"),
   509 => (x"5b",x"5e",x"0e",x"87"),
   510 => (x"f8",x"0e",x"5d",x"5c"),
   511 => (x"9c",x"4c",x"71",x"86"),
   512 => (x"c0",x"87",x"c5",x"05"),
   513 => (x"87",x"c0",x"c3",x"48"),
   514 => (x"48",x"7e",x"a4",x"c8"),
   515 => (x"66",x"d8",x"78",x"c0"),
   516 => (x"d8",x"87",x"c7",x"02"),
   517 => (x"05",x"bf",x"97",x"66"),
   518 => (x"48",x"c0",x"87",x"c5"),
   519 => (x"c0",x"87",x"e9",x"c2"),
   520 => (x"49",x"49",x"c1",x"1e"),
   521 => (x"c4",x"87",x"d3",x"ca"),
   522 => (x"9d",x"4d",x"70",x"86"),
   523 => (x"87",x"c2",x"c1",x"02"),
   524 => (x"4a",x"d6",x"e3",x"c2"),
   525 => (x"e0",x"49",x"66",x"d8"),
   526 => (x"98",x"70",x"87",x"d4"),
   527 => (x"87",x"f2",x"c0",x"02"),
   528 => (x"66",x"d8",x"4a",x"75"),
   529 => (x"e0",x"4b",x"cb",x"49"),
   530 => (x"98",x"70",x"87",x"f9"),
   531 => (x"87",x"e2",x"c0",x"02"),
   532 => (x"9d",x"75",x"1e",x"c0"),
   533 => (x"c8",x"87",x"c7",x"02"),
   534 => (x"78",x"c0",x"48",x"a6"),
   535 => (x"a6",x"c8",x"87",x"c5"),
   536 => (x"c8",x"78",x"c1",x"48"),
   537 => (x"d1",x"c9",x"49",x"66"),
   538 => (x"70",x"86",x"c4",x"87"),
   539 => (x"fe",x"05",x"9d",x"4d"),
   540 => (x"9d",x"75",x"87",x"fe"),
   541 => (x"87",x"ce",x"c1",x"02"),
   542 => (x"6e",x"49",x"a5",x"dc"),
   543 => (x"da",x"78",x"69",x"48"),
   544 => (x"a6",x"c4",x"49",x"a5"),
   545 => (x"78",x"a4",x"c4",x"48"),
   546 => (x"c4",x"48",x"69",x"9f"),
   547 => (x"c2",x"78",x"08",x"66"),
   548 => (x"02",x"bf",x"ce",x"e3"),
   549 => (x"a5",x"d4",x"87",x"d2"),
   550 => (x"49",x"69",x"9f",x"49"),
   551 => (x"99",x"ff",x"ff",x"c0"),
   552 => (x"30",x"d0",x"48",x"71"),
   553 => (x"87",x"c2",x"7e",x"70"),
   554 => (x"48",x"6e",x"7e",x"c0"),
   555 => (x"80",x"bf",x"66",x"c4"),
   556 => (x"78",x"08",x"66",x"c4"),
   557 => (x"a4",x"cc",x"7c",x"c0"),
   558 => (x"bf",x"66",x"c4",x"49"),
   559 => (x"49",x"a4",x"d0",x"79"),
   560 => (x"48",x"c1",x"79",x"c0"),
   561 => (x"48",x"c0",x"87",x"c2"),
   562 => (x"ee",x"fa",x"8e",x"f8"),
   563 => (x"5b",x"5e",x"0e",x"87"),
   564 => (x"4c",x"71",x"0e",x"5c"),
   565 => (x"cb",x"c1",x"02",x"9c"),
   566 => (x"49",x"a4",x"c8",x"87"),
   567 => (x"c3",x"c1",x"02",x"69"),
   568 => (x"cc",x"49",x"6c",x"87"),
   569 => (x"80",x"71",x"48",x"66"),
   570 => (x"70",x"58",x"a6",x"d0"),
   571 => (x"ca",x"e3",x"c2",x"b9"),
   572 => (x"ba",x"ff",x"4a",x"bf"),
   573 => (x"99",x"71",x"99",x"72"),
   574 => (x"87",x"e5",x"c0",x"02"),
   575 => (x"6b",x"4b",x"a4",x"c4"),
   576 => (x"87",x"ff",x"f9",x"49"),
   577 => (x"e3",x"c2",x"7b",x"70"),
   578 => (x"6c",x"49",x"bf",x"c6"),
   579 => (x"cc",x"7c",x"71",x"81"),
   580 => (x"e3",x"c2",x"b9",x"66"),
   581 => (x"ff",x"4a",x"bf",x"ca"),
   582 => (x"71",x"99",x"72",x"ba"),
   583 => (x"db",x"ff",x"05",x"99"),
   584 => (x"7c",x"66",x"cc",x"87"),
   585 => (x"1e",x"87",x"d6",x"f9"),
   586 => (x"4b",x"71",x"1e",x"73"),
   587 => (x"87",x"c7",x"02",x"9b"),
   588 => (x"69",x"49",x"a3",x"c8"),
   589 => (x"c0",x"87",x"c5",x"05"),
   590 => (x"87",x"f6",x"c0",x"48"),
   591 => (x"bf",x"df",x"e7",x"c2"),
   592 => (x"4a",x"a3",x"c4",x"49"),
   593 => (x"8a",x"c2",x"4a",x"6a"),
   594 => (x"bf",x"c6",x"e3",x"c2"),
   595 => (x"49",x"a1",x"72",x"92"),
   596 => (x"bf",x"ca",x"e3",x"c2"),
   597 => (x"72",x"9a",x"6b",x"4a"),
   598 => (x"f2",x"c0",x"49",x"a1"),
   599 => (x"66",x"c8",x"59",x"d5"),
   600 => (x"e6",x"ea",x"71",x"1e"),
   601 => (x"70",x"86",x"c4",x"87"),
   602 => (x"87",x"c4",x"05",x"98"),
   603 => (x"87",x"c2",x"48",x"c0"),
   604 => (x"ca",x"f8",x"48",x"c1"),
   605 => (x"1e",x"73",x"1e",x"87"),
   606 => (x"02",x"9b",x"4b",x"71"),
   607 => (x"a3",x"c8",x"87",x"c7"),
   608 => (x"c5",x"05",x"69",x"49"),
   609 => (x"c0",x"48",x"c0",x"87"),
   610 => (x"e7",x"c2",x"87",x"f6"),
   611 => (x"c4",x"49",x"bf",x"df"),
   612 => (x"4a",x"6a",x"4a",x"a3"),
   613 => (x"e3",x"c2",x"8a",x"c2"),
   614 => (x"72",x"92",x"bf",x"c6"),
   615 => (x"e3",x"c2",x"49",x"a1"),
   616 => (x"6b",x"4a",x"bf",x"ca"),
   617 => (x"49",x"a1",x"72",x"9a"),
   618 => (x"59",x"d5",x"f2",x"c0"),
   619 => (x"71",x"1e",x"66",x"c8"),
   620 => (x"c4",x"87",x"d1",x"e6"),
   621 => (x"05",x"98",x"70",x"86"),
   622 => (x"48",x"c0",x"87",x"c4"),
   623 => (x"48",x"c1",x"87",x"c2"),
   624 => (x"0e",x"87",x"fc",x"f6"),
   625 => (x"5d",x"5c",x"5b",x"5e"),
   626 => (x"4b",x"71",x"1e",x"0e"),
   627 => (x"73",x"4d",x"66",x"d4"),
   628 => (x"cc",x"c1",x"02",x"9b"),
   629 => (x"49",x"a3",x"c8",x"87"),
   630 => (x"c4",x"c1",x"02",x"69"),
   631 => (x"4c",x"a3",x"d0",x"87"),
   632 => (x"bf",x"ca",x"e3",x"c2"),
   633 => (x"6c",x"b9",x"ff",x"49"),
   634 => (x"d4",x"7e",x"99",x"4a"),
   635 => (x"cd",x"06",x"a9",x"66"),
   636 => (x"7c",x"7b",x"c0",x"87"),
   637 => (x"c4",x"4a",x"a3",x"cc"),
   638 => (x"79",x"6a",x"49",x"a3"),
   639 => (x"49",x"72",x"87",x"ca"),
   640 => (x"d4",x"99",x"c0",x"f8"),
   641 => (x"8d",x"71",x"4d",x"66"),
   642 => (x"29",x"c9",x"49",x"75"),
   643 => (x"49",x"73",x"1e",x"71"),
   644 => (x"c2",x"87",x"fa",x"fa"),
   645 => (x"73",x"1e",x"c6",x"db"),
   646 => (x"87",x"cb",x"fc",x"49"),
   647 => (x"66",x"d4",x"86",x"c8"),
   648 => (x"d6",x"f5",x"26",x"7c"),
   649 => (x"1e",x"73",x"1e",x"87"),
   650 => (x"02",x"9b",x"4b",x"71"),
   651 => (x"c2",x"87",x"e4",x"c0"),
   652 => (x"73",x"5b",x"f3",x"e7"),
   653 => (x"c2",x"8a",x"c2",x"4a"),
   654 => (x"49",x"bf",x"c6",x"e3"),
   655 => (x"df",x"e7",x"c2",x"92"),
   656 => (x"80",x"72",x"48",x"bf"),
   657 => (x"58",x"f7",x"e7",x"c2"),
   658 => (x"30",x"c4",x"48",x"71"),
   659 => (x"58",x"d6",x"e3",x"c2"),
   660 => (x"c2",x"87",x"ed",x"c0"),
   661 => (x"c2",x"48",x"ef",x"e7"),
   662 => (x"78",x"bf",x"e3",x"e7"),
   663 => (x"48",x"f3",x"e7",x"c2"),
   664 => (x"bf",x"e7",x"e7",x"c2"),
   665 => (x"ce",x"e3",x"c2",x"78"),
   666 => (x"87",x"c9",x"02",x"bf"),
   667 => (x"bf",x"c6",x"e3",x"c2"),
   668 => (x"c7",x"31",x"c4",x"49"),
   669 => (x"eb",x"e7",x"c2",x"87"),
   670 => (x"31",x"c4",x"49",x"bf"),
   671 => (x"59",x"d6",x"e3",x"c2"),
   672 => (x"0e",x"87",x"fc",x"f3"),
   673 => (x"0e",x"5c",x"5b",x"5e"),
   674 => (x"4b",x"c0",x"4a",x"71"),
   675 => (x"c0",x"02",x"9a",x"72"),
   676 => (x"a2",x"da",x"87",x"e0"),
   677 => (x"4b",x"69",x"9f",x"49"),
   678 => (x"bf",x"ce",x"e3",x"c2"),
   679 => (x"d4",x"87",x"cf",x"02"),
   680 => (x"69",x"9f",x"49",x"a2"),
   681 => (x"ff",x"c0",x"4c",x"49"),
   682 => (x"34",x"d0",x"9c",x"ff"),
   683 => (x"4c",x"c0",x"87",x"c2"),
   684 => (x"49",x"73",x"b3",x"74"),
   685 => (x"f3",x"87",x"ee",x"fd"),
   686 => (x"5e",x"0e",x"87",x"c3"),
   687 => (x"0e",x"5d",x"5c",x"5b"),
   688 => (x"4a",x"71",x"86",x"f4"),
   689 => (x"9a",x"72",x"7e",x"c0"),
   690 => (x"c2",x"87",x"d8",x"02"),
   691 => (x"c0",x"48",x"c2",x"db"),
   692 => (x"fa",x"da",x"c2",x"78"),
   693 => (x"f3",x"e7",x"c2",x"48"),
   694 => (x"da",x"c2",x"78",x"bf"),
   695 => (x"e7",x"c2",x"48",x"fe"),
   696 => (x"c2",x"78",x"bf",x"ef"),
   697 => (x"c0",x"48",x"e3",x"e3"),
   698 => (x"d2",x"e3",x"c2",x"50"),
   699 => (x"db",x"c2",x"49",x"bf"),
   700 => (x"71",x"4a",x"bf",x"c2"),
   701 => (x"c9",x"c4",x"03",x"aa"),
   702 => (x"cf",x"49",x"72",x"87"),
   703 => (x"e9",x"c0",x"05",x"99"),
   704 => (x"d1",x"f2",x"c0",x"87"),
   705 => (x"fa",x"da",x"c2",x"48"),
   706 => (x"db",x"c2",x"78",x"bf"),
   707 => (x"da",x"c2",x"1e",x"c6"),
   708 => (x"c2",x"49",x"bf",x"fa"),
   709 => (x"c1",x"48",x"fa",x"da"),
   710 => (x"e3",x"71",x"78",x"a1"),
   711 => (x"86",x"c4",x"87",x"ed"),
   712 => (x"48",x"cd",x"f2",x"c0"),
   713 => (x"78",x"c6",x"db",x"c2"),
   714 => (x"f2",x"c0",x"87",x"cc"),
   715 => (x"c0",x"48",x"bf",x"cd"),
   716 => (x"f2",x"c0",x"80",x"e0"),
   717 => (x"db",x"c2",x"58",x"d1"),
   718 => (x"c1",x"48",x"bf",x"c2"),
   719 => (x"c6",x"db",x"c2",x"80"),
   720 => (x"0c",x"8d",x"27",x"58"),
   721 => (x"97",x"bf",x"00",x"00"),
   722 => (x"02",x"9d",x"4d",x"bf"),
   723 => (x"c3",x"87",x"e3",x"c2"),
   724 => (x"c2",x"02",x"ad",x"e5"),
   725 => (x"f2",x"c0",x"87",x"dc"),
   726 => (x"cb",x"4b",x"bf",x"cd"),
   727 => (x"4c",x"11",x"49",x"a3"),
   728 => (x"c1",x"05",x"ac",x"cf"),
   729 => (x"49",x"75",x"87",x"d2"),
   730 => (x"89",x"c1",x"99",x"df"),
   731 => (x"e3",x"c2",x"91",x"cd"),
   732 => (x"a3",x"c1",x"81",x"d6"),
   733 => (x"c3",x"51",x"12",x"4a"),
   734 => (x"51",x"12",x"4a",x"a3"),
   735 => (x"12",x"4a",x"a3",x"c5"),
   736 => (x"4a",x"a3",x"c7",x"51"),
   737 => (x"a3",x"c9",x"51",x"12"),
   738 => (x"ce",x"51",x"12",x"4a"),
   739 => (x"51",x"12",x"4a",x"a3"),
   740 => (x"12",x"4a",x"a3",x"d0"),
   741 => (x"4a",x"a3",x"d2",x"51"),
   742 => (x"a3",x"d4",x"51",x"12"),
   743 => (x"d6",x"51",x"12",x"4a"),
   744 => (x"51",x"12",x"4a",x"a3"),
   745 => (x"12",x"4a",x"a3",x"d8"),
   746 => (x"4a",x"a3",x"dc",x"51"),
   747 => (x"a3",x"de",x"51",x"12"),
   748 => (x"c1",x"51",x"12",x"4a"),
   749 => (x"87",x"fa",x"c0",x"7e"),
   750 => (x"99",x"c8",x"49",x"74"),
   751 => (x"87",x"eb",x"c0",x"05"),
   752 => (x"99",x"d0",x"49",x"74"),
   753 => (x"dc",x"87",x"d1",x"05"),
   754 => (x"cb",x"c0",x"02",x"66"),
   755 => (x"dc",x"49",x"73",x"87"),
   756 => (x"98",x"70",x"0f",x"66"),
   757 => (x"87",x"d3",x"c0",x"02"),
   758 => (x"c6",x"c0",x"05",x"6e"),
   759 => (x"d6",x"e3",x"c2",x"87"),
   760 => (x"c0",x"50",x"c0",x"48"),
   761 => (x"48",x"bf",x"cd",x"f2"),
   762 => (x"c2",x"87",x"dd",x"c2"),
   763 => (x"c0",x"48",x"e3",x"e3"),
   764 => (x"e3",x"c2",x"7e",x"50"),
   765 => (x"c2",x"49",x"bf",x"d2"),
   766 => (x"4a",x"bf",x"c2",x"db"),
   767 => (x"fb",x"04",x"aa",x"71"),
   768 => (x"e7",x"c2",x"87",x"f7"),
   769 => (x"c0",x"05",x"bf",x"f3"),
   770 => (x"e3",x"c2",x"87",x"c8"),
   771 => (x"c1",x"02",x"bf",x"ce"),
   772 => (x"da",x"c2",x"87",x"f4"),
   773 => (x"ed",x"49",x"bf",x"fe"),
   774 => (x"db",x"c2",x"87",x"e9"),
   775 => (x"a6",x"c4",x"58",x"c2"),
   776 => (x"fe",x"da",x"c2",x"48"),
   777 => (x"e3",x"c2",x"78",x"bf"),
   778 => (x"c0",x"02",x"bf",x"ce"),
   779 => (x"66",x"c4",x"87",x"d8"),
   780 => (x"ff",x"ff",x"cf",x"49"),
   781 => (x"a9",x"99",x"f8",x"ff"),
   782 => (x"87",x"c5",x"c0",x"02"),
   783 => (x"e1",x"c0",x"4c",x"c0"),
   784 => (x"c0",x"4c",x"c1",x"87"),
   785 => (x"66",x"c4",x"87",x"dc"),
   786 => (x"f8",x"ff",x"cf",x"49"),
   787 => (x"c0",x"02",x"a9",x"99"),
   788 => (x"a6",x"c8",x"87",x"c8"),
   789 => (x"c0",x"78",x"c0",x"48"),
   790 => (x"a6",x"c8",x"87",x"c5"),
   791 => (x"c8",x"78",x"c1",x"48"),
   792 => (x"9c",x"74",x"4c",x"66"),
   793 => (x"87",x"de",x"c0",x"05"),
   794 => (x"c2",x"49",x"66",x"c4"),
   795 => (x"c6",x"e3",x"c2",x"89"),
   796 => (x"e7",x"c2",x"91",x"bf"),
   797 => (x"71",x"48",x"bf",x"df"),
   798 => (x"fe",x"da",x"c2",x"80"),
   799 => (x"c2",x"db",x"c2",x"58"),
   800 => (x"f9",x"78",x"c0",x"48"),
   801 => (x"48",x"c0",x"87",x"e3"),
   802 => (x"ee",x"eb",x"8e",x"f4"),
   803 => (x"00",x"00",x"00",x"87"),
   804 => (x"ff",x"ff",x"ff",x"00"),
   805 => (x"00",x"0c",x"9d",x"ff"),
   806 => (x"00",x"0c",x"a6",x"00"),
   807 => (x"54",x"41",x"46",x"00"),
   808 => (x"20",x"20",x"32",x"33"),
   809 => (x"41",x"46",x"00",x"20"),
   810 => (x"20",x"36",x"31",x"54"),
   811 => (x"1e",x"00",x"20",x"20"),
   812 => (x"c3",x"48",x"d4",x"ff"),
   813 => (x"48",x"68",x"78",x"ff"),
   814 => (x"ff",x"1e",x"4f",x"26"),
   815 => (x"ff",x"c3",x"48",x"d4"),
   816 => (x"48",x"d0",x"ff",x"78"),
   817 => (x"ff",x"78",x"e1",x"c0"),
   818 => (x"78",x"d4",x"48",x"d4"),
   819 => (x"48",x"f7",x"e7",x"c2"),
   820 => (x"50",x"bf",x"d4",x"ff"),
   821 => (x"ff",x"1e",x"4f",x"26"),
   822 => (x"e0",x"c0",x"48",x"d0"),
   823 => (x"1e",x"4f",x"26",x"78"),
   824 => (x"70",x"87",x"cc",x"ff"),
   825 => (x"c6",x"02",x"99",x"49"),
   826 => (x"a9",x"fb",x"c0",x"87"),
   827 => (x"71",x"87",x"f1",x"05"),
   828 => (x"0e",x"4f",x"26",x"48"),
   829 => (x"0e",x"5c",x"5b",x"5e"),
   830 => (x"4c",x"c0",x"4b",x"71"),
   831 => (x"70",x"87",x"f0",x"fe"),
   832 => (x"c0",x"02",x"99",x"49"),
   833 => (x"ec",x"c0",x"87",x"f9"),
   834 => (x"f2",x"c0",x"02",x"a9"),
   835 => (x"a9",x"fb",x"c0",x"87"),
   836 => (x"87",x"eb",x"c0",x"02"),
   837 => (x"ac",x"b7",x"66",x"cc"),
   838 => (x"d0",x"87",x"c7",x"03"),
   839 => (x"87",x"c2",x"02",x"66"),
   840 => (x"99",x"71",x"53",x"71"),
   841 => (x"c1",x"87",x"c2",x"02"),
   842 => (x"87",x"c3",x"fe",x"84"),
   843 => (x"02",x"99",x"49",x"70"),
   844 => (x"ec",x"c0",x"87",x"cd"),
   845 => (x"87",x"c7",x"02",x"a9"),
   846 => (x"05",x"a9",x"fb",x"c0"),
   847 => (x"d0",x"87",x"d5",x"ff"),
   848 => (x"87",x"c3",x"02",x"66"),
   849 => (x"c0",x"7b",x"97",x"c0"),
   850 => (x"c4",x"05",x"a9",x"ec"),
   851 => (x"c5",x"4a",x"74",x"87"),
   852 => (x"c0",x"4a",x"74",x"87"),
   853 => (x"48",x"72",x"8a",x"0a"),
   854 => (x"4d",x"26",x"87",x"c2"),
   855 => (x"4b",x"26",x"4c",x"26"),
   856 => (x"fd",x"1e",x"4f",x"26"),
   857 => (x"49",x"70",x"87",x"c9"),
   858 => (x"aa",x"f0",x"c0",x"4a"),
   859 => (x"c0",x"87",x"c9",x"04"),
   860 => (x"c3",x"01",x"aa",x"f9"),
   861 => (x"8a",x"f0",x"c0",x"87"),
   862 => (x"04",x"aa",x"c1",x"c1"),
   863 => (x"da",x"c1",x"87",x"c9"),
   864 => (x"87",x"c3",x"01",x"aa"),
   865 => (x"72",x"8a",x"f7",x"c0"),
   866 => (x"0e",x"4f",x"26",x"48"),
   867 => (x"5d",x"5c",x"5b",x"5e"),
   868 => (x"71",x"86",x"f8",x"0e"),
   869 => (x"fc",x"4d",x"c0",x"4c"),
   870 => (x"4b",x"c0",x"87",x"e0"),
   871 => (x"97",x"ea",x"f8",x"c0"),
   872 => (x"a9",x"c0",x"49",x"bf"),
   873 => (x"fc",x"87",x"cf",x"04"),
   874 => (x"83",x"c1",x"87",x"f5"),
   875 => (x"97",x"ea",x"f8",x"c0"),
   876 => (x"06",x"ab",x"49",x"bf"),
   877 => (x"f8",x"c0",x"87",x"f1"),
   878 => (x"02",x"bf",x"97",x"ea"),
   879 => (x"ee",x"fb",x"87",x"cf"),
   880 => (x"99",x"49",x"70",x"87"),
   881 => (x"c0",x"87",x"c6",x"02"),
   882 => (x"f1",x"05",x"a9",x"ec"),
   883 => (x"fb",x"4b",x"c0",x"87"),
   884 => (x"7e",x"70",x"87",x"dd"),
   885 => (x"c8",x"87",x"d8",x"fb"),
   886 => (x"d2",x"fb",x"58",x"a6"),
   887 => (x"c1",x"4a",x"70",x"87"),
   888 => (x"49",x"a4",x"c8",x"83"),
   889 => (x"6e",x"49",x"69",x"97"),
   890 => (x"87",x"da",x"05",x"a9"),
   891 => (x"97",x"49",x"a4",x"c9"),
   892 => (x"66",x"c4",x"49",x"69"),
   893 => (x"87",x"ce",x"05",x"a9"),
   894 => (x"97",x"49",x"a4",x"ca"),
   895 => (x"05",x"aa",x"49",x"69"),
   896 => (x"4d",x"c1",x"87",x"c4"),
   897 => (x"48",x"6e",x"87",x"d4"),
   898 => (x"02",x"a8",x"ec",x"c0"),
   899 => (x"48",x"6e",x"87",x"c8"),
   900 => (x"05",x"a8",x"fb",x"c0"),
   901 => (x"4b",x"c0",x"87",x"c4"),
   902 => (x"9d",x"75",x"4d",x"c1"),
   903 => (x"87",x"ef",x"fe",x"02"),
   904 => (x"73",x"87",x"f3",x"fa"),
   905 => (x"fc",x"8e",x"f8",x"48"),
   906 => (x"0e",x"00",x"87",x"f0"),
   907 => (x"5d",x"5c",x"5b",x"5e"),
   908 => (x"71",x"86",x"f8",x"0e"),
   909 => (x"4b",x"d4",x"ff",x"7e"),
   910 => (x"e7",x"c2",x"1e",x"6e"),
   911 => (x"f4",x"e6",x"49",x"fc"),
   912 => (x"70",x"86",x"c4",x"87"),
   913 => (x"ea",x"c4",x"02",x"98"),
   914 => (x"da",x"e3",x"c1",x"87"),
   915 => (x"49",x"6e",x"4d",x"bf"),
   916 => (x"c8",x"87",x"f8",x"fc"),
   917 => (x"98",x"70",x"58",x"a6"),
   918 => (x"c4",x"87",x"c5",x"05"),
   919 => (x"78",x"c1",x"48",x"a6"),
   920 => (x"c5",x"48",x"d0",x"ff"),
   921 => (x"7b",x"d5",x"c1",x"78"),
   922 => (x"c1",x"49",x"66",x"c4"),
   923 => (x"c1",x"31",x"c6",x"89"),
   924 => (x"bf",x"97",x"d8",x"e3"),
   925 => (x"b0",x"71",x"48",x"4a"),
   926 => (x"d0",x"ff",x"7b",x"70"),
   927 => (x"c2",x"78",x"c4",x"48"),
   928 => (x"bf",x"97",x"f7",x"e7"),
   929 => (x"02",x"99",x"d0",x"49"),
   930 => (x"78",x"c5",x"87",x"d7"),
   931 => (x"c0",x"7b",x"d6",x"c1"),
   932 => (x"7b",x"ff",x"c3",x"4a"),
   933 => (x"e0",x"c0",x"82",x"c1"),
   934 => (x"87",x"f5",x"04",x"aa"),
   935 => (x"c4",x"48",x"d0",x"ff"),
   936 => (x"7b",x"ff",x"c3",x"78"),
   937 => (x"c5",x"48",x"d0",x"ff"),
   938 => (x"7b",x"d3",x"c1",x"78"),
   939 => (x"78",x"c4",x"7b",x"c1"),
   940 => (x"06",x"ad",x"b7",x"c0"),
   941 => (x"c2",x"87",x"eb",x"c2"),
   942 => (x"4c",x"bf",x"c4",x"e8"),
   943 => (x"c2",x"02",x"9c",x"8d"),
   944 => (x"db",x"c2",x"87",x"c2"),
   945 => (x"a6",x"c4",x"7e",x"c6"),
   946 => (x"78",x"c0",x"c8",x"48"),
   947 => (x"ac",x"b7",x"c0",x"8c"),
   948 => (x"c8",x"87",x"c6",x"03"),
   949 => (x"c0",x"78",x"a4",x"c0"),
   950 => (x"f7",x"e7",x"c2",x"4c"),
   951 => (x"d0",x"49",x"bf",x"97"),
   952 => (x"87",x"d0",x"02",x"99"),
   953 => (x"e7",x"c2",x"1e",x"c0"),
   954 => (x"fa",x"e8",x"49",x"fc"),
   955 => (x"70",x"86",x"c4",x"87"),
   956 => (x"87",x"f5",x"c0",x"4a"),
   957 => (x"1e",x"c6",x"db",x"c2"),
   958 => (x"49",x"fc",x"e7",x"c2"),
   959 => (x"c4",x"87",x"e8",x"e8"),
   960 => (x"ff",x"4a",x"70",x"86"),
   961 => (x"c5",x"c8",x"48",x"d0"),
   962 => (x"7b",x"d4",x"c1",x"78"),
   963 => (x"7b",x"bf",x"97",x"6e"),
   964 => (x"80",x"c1",x"48",x"6e"),
   965 => (x"66",x"c4",x"7e",x"70"),
   966 => (x"c8",x"88",x"c1",x"48"),
   967 => (x"98",x"70",x"58",x"a6"),
   968 => (x"87",x"e8",x"ff",x"05"),
   969 => (x"c4",x"48",x"d0",x"ff"),
   970 => (x"05",x"9a",x"72",x"78"),
   971 => (x"48",x"c0",x"87",x"c5"),
   972 => (x"c1",x"87",x"c2",x"c1"),
   973 => (x"fc",x"e7",x"c2",x"1e"),
   974 => (x"87",x"d1",x"e6",x"49"),
   975 => (x"9c",x"74",x"86",x"c4"),
   976 => (x"87",x"fe",x"fd",x"05"),
   977 => (x"06",x"ad",x"b7",x"c0"),
   978 => (x"e7",x"c2",x"87",x"d1"),
   979 => (x"78",x"c0",x"48",x"fc"),
   980 => (x"78",x"c0",x"80",x"d0"),
   981 => (x"e8",x"c2",x"80",x"f4"),
   982 => (x"c0",x"78",x"bf",x"c8"),
   983 => (x"fd",x"01",x"ad",x"b7"),
   984 => (x"d0",x"ff",x"87",x"d5"),
   985 => (x"c1",x"78",x"c5",x"48"),
   986 => (x"7b",x"c0",x"7b",x"d3"),
   987 => (x"48",x"c1",x"78",x"c4"),
   988 => (x"c0",x"87",x"c2",x"c0"),
   989 => (x"26",x"8e",x"f8",x"48"),
   990 => (x"26",x"4c",x"26",x"4d"),
   991 => (x"0e",x"4f",x"26",x"4b"),
   992 => (x"5d",x"5c",x"5b",x"5e"),
   993 => (x"4b",x"71",x"1e",x"0e"),
   994 => (x"ab",x"4d",x"4c",x"c0"),
   995 => (x"87",x"e8",x"c0",x"04"),
   996 => (x"1e",x"cb",x"f6",x"c0"),
   997 => (x"c4",x"02",x"9d",x"75"),
   998 => (x"c2",x"4a",x"c0",x"87"),
   999 => (x"72",x"4a",x"c1",x"87"),
  1000 => (x"87",x"d6",x"ec",x"49"),
  1001 => (x"7e",x"70",x"86",x"c4"),
  1002 => (x"05",x"6e",x"84",x"c1"),
  1003 => (x"4c",x"73",x"87",x"c2"),
  1004 => (x"ac",x"73",x"85",x"c1"),
  1005 => (x"87",x"d8",x"ff",x"06"),
  1006 => (x"fe",x"26",x"48",x"6e"),
  1007 => (x"5e",x"0e",x"87",x"f9"),
  1008 => (x"71",x"0e",x"5c",x"5b"),
  1009 => (x"02",x"66",x"cc",x"4b"),
  1010 => (x"c0",x"4c",x"87",x"d8"),
  1011 => (x"d8",x"02",x"8c",x"f0"),
  1012 => (x"c1",x"4a",x"74",x"87"),
  1013 => (x"87",x"d1",x"02",x"8a"),
  1014 => (x"87",x"cd",x"02",x"8a"),
  1015 => (x"87",x"c9",x"02",x"8a"),
  1016 => (x"49",x"73",x"87",x"d9"),
  1017 => (x"d2",x"87",x"c4",x"f9"),
  1018 => (x"c0",x"1e",x"74",x"87"),
  1019 => (x"f7",x"d8",x"c1",x"49"),
  1020 => (x"73",x"1e",x"74",x"87"),
  1021 => (x"ef",x"d8",x"c1",x"49"),
  1022 => (x"fd",x"86",x"c8",x"87"),
  1023 => (x"5e",x"0e",x"87",x"fb"),
  1024 => (x"0e",x"5d",x"5c",x"5b"),
  1025 => (x"49",x"4c",x"71",x"1e"),
  1026 => (x"e8",x"c2",x"91",x"de"),
  1027 => (x"85",x"71",x"4d",x"e4"),
  1028 => (x"c1",x"02",x"6d",x"97"),
  1029 => (x"e8",x"c2",x"87",x"dc"),
  1030 => (x"74",x"49",x"bf",x"d0"),
  1031 => (x"de",x"fd",x"71",x"81"),
  1032 => (x"48",x"7e",x"70",x"87"),
  1033 => (x"f2",x"c0",x"02",x"98"),
  1034 => (x"d8",x"e8",x"c2",x"87"),
  1035 => (x"cb",x"4a",x"70",x"4b"),
  1036 => (x"f2",x"c1",x"ff",x"49"),
  1037 => (x"cb",x"4b",x"74",x"87"),
  1038 => (x"ec",x"e3",x"c1",x"93"),
  1039 => (x"c1",x"83",x"c4",x"83"),
  1040 => (x"74",x"7b",x"f6",x"c1"),
  1041 => (x"d0",x"c1",x"c1",x"49"),
  1042 => (x"c1",x"7b",x"75",x"87"),
  1043 => (x"bf",x"97",x"d9",x"e3"),
  1044 => (x"e8",x"c2",x"1e",x"49"),
  1045 => (x"e5",x"fd",x"49",x"d8"),
  1046 => (x"74",x"86",x"c4",x"87"),
  1047 => (x"f8",x"c0",x"c1",x"49"),
  1048 => (x"c1",x"49",x"c0",x"87"),
  1049 => (x"c2",x"87",x"d7",x"c2"),
  1050 => (x"c0",x"48",x"f8",x"e7"),
  1051 => (x"de",x"49",x"c1",x"78"),
  1052 => (x"fc",x"26",x"87",x"cd"),
  1053 => (x"6f",x"4c",x"87",x"c1"),
  1054 => (x"6e",x"69",x"64",x"61"),
  1055 => (x"2e",x"2e",x"2e",x"67"),
  1056 => (x"1e",x"73",x"1e",x"00"),
  1057 => (x"c2",x"49",x"4a",x"71"),
  1058 => (x"81",x"bf",x"d0",x"e8"),
  1059 => (x"87",x"ef",x"fb",x"71"),
  1060 => (x"02",x"9b",x"4b",x"70"),
  1061 => (x"e7",x"49",x"87",x"c4"),
  1062 => (x"e8",x"c2",x"87",x"e9"),
  1063 => (x"78",x"c0",x"48",x"d0"),
  1064 => (x"da",x"dd",x"49",x"c1"),
  1065 => (x"87",x"d3",x"fb",x"87"),
  1066 => (x"c1",x"49",x"c0",x"1e"),
  1067 => (x"26",x"87",x"cf",x"c1"),
  1068 => (x"4a",x"71",x"1e",x"4f"),
  1069 => (x"c1",x"91",x"cb",x"49"),
  1070 => (x"c8",x"81",x"ec",x"e3"),
  1071 => (x"c2",x"48",x"11",x"81"),
  1072 => (x"c2",x"58",x"fc",x"e7"),
  1073 => (x"c0",x"48",x"d0",x"e8"),
  1074 => (x"dc",x"49",x"c1",x"78"),
  1075 => (x"4f",x"26",x"87",x"f1"),
  1076 => (x"02",x"99",x"71",x"1e"),
  1077 => (x"e5",x"c1",x"87",x"d2"),
  1078 => (x"50",x"c0",x"48",x"c1"),
  1079 => (x"c2",x"c1",x"80",x"f7"),
  1080 => (x"e3",x"c1",x"40",x"f1"),
  1081 => (x"87",x"ce",x"78",x"e5"),
  1082 => (x"48",x"fd",x"e4",x"c1"),
  1083 => (x"78",x"de",x"e3",x"c1"),
  1084 => (x"c2",x"c1",x"80",x"fc"),
  1085 => (x"4f",x"26",x"78",x"e8"),
  1086 => (x"5c",x"5b",x"5e",x"0e"),
  1087 => (x"86",x"f4",x"0e",x"5d"),
  1088 => (x"4d",x"c6",x"db",x"c2"),
  1089 => (x"a6",x"c4",x"4c",x"c0"),
  1090 => (x"c2",x"78",x"c0",x"48"),
  1091 => (x"48",x"bf",x"d0",x"e8"),
  1092 => (x"c1",x"06",x"a8",x"c0"),
  1093 => (x"db",x"c2",x"87",x"c0"),
  1094 => (x"02",x"98",x"48",x"c6"),
  1095 => (x"c0",x"87",x"f7",x"c0"),
  1096 => (x"c8",x"1e",x"cb",x"f6"),
  1097 => (x"87",x"c7",x"02",x"66"),
  1098 => (x"c0",x"48",x"a6",x"c4"),
  1099 => (x"c4",x"87",x"c5",x"78"),
  1100 => (x"78",x"c1",x"48",x"a6"),
  1101 => (x"e6",x"49",x"66",x"c4"),
  1102 => (x"86",x"c4",x"87",x"c0"),
  1103 => (x"84",x"c1",x"4d",x"70"),
  1104 => (x"c1",x"48",x"66",x"c4"),
  1105 => (x"58",x"a6",x"c8",x"80"),
  1106 => (x"bf",x"d0",x"e8",x"c2"),
  1107 => (x"87",x"c6",x"03",x"ac"),
  1108 => (x"ff",x"05",x"9d",x"75"),
  1109 => (x"4c",x"c0",x"87",x"c9"),
  1110 => (x"c3",x"02",x"9d",x"75"),
  1111 => (x"f6",x"c0",x"87",x"dc"),
  1112 => (x"66",x"c8",x"1e",x"cb"),
  1113 => (x"cc",x"87",x"c7",x"02"),
  1114 => (x"78",x"c0",x"48",x"a6"),
  1115 => (x"a6",x"cc",x"87",x"c5"),
  1116 => (x"cc",x"78",x"c1",x"48"),
  1117 => (x"c1",x"e5",x"49",x"66"),
  1118 => (x"70",x"86",x"c4",x"87"),
  1119 => (x"02",x"98",x"48",x"7e"),
  1120 => (x"49",x"87",x"e4",x"c2"),
  1121 => (x"69",x"97",x"81",x"cb"),
  1122 => (x"02",x"99",x"d0",x"49"),
  1123 => (x"74",x"87",x"d4",x"c1"),
  1124 => (x"c1",x"91",x"cb",x"49"),
  1125 => (x"c1",x"81",x"ec",x"e3"),
  1126 => (x"c8",x"79",x"c1",x"c2"),
  1127 => (x"51",x"ff",x"c3",x"81"),
  1128 => (x"91",x"de",x"49",x"74"),
  1129 => (x"4d",x"e4",x"e8",x"c2"),
  1130 => (x"c1",x"c2",x"85",x"71"),
  1131 => (x"a5",x"c1",x"7d",x"97"),
  1132 => (x"51",x"e0",x"c0",x"49"),
  1133 => (x"97",x"d6",x"e3",x"c2"),
  1134 => (x"87",x"d2",x"02",x"bf"),
  1135 => (x"a5",x"c2",x"84",x"c1"),
  1136 => (x"d6",x"e3",x"c2",x"4b"),
  1137 => (x"fe",x"49",x"db",x"4a"),
  1138 => (x"c1",x"87",x"dc",x"fb"),
  1139 => (x"a5",x"cd",x"87",x"d9"),
  1140 => (x"c1",x"51",x"c0",x"49"),
  1141 => (x"4b",x"a5",x"c2",x"84"),
  1142 => (x"49",x"cb",x"4a",x"6e"),
  1143 => (x"87",x"c7",x"fb",x"fe"),
  1144 => (x"74",x"87",x"c4",x"c1"),
  1145 => (x"c1",x"91",x"cb",x"49"),
  1146 => (x"c0",x"81",x"ec",x"e3"),
  1147 => (x"c2",x"79",x"fe",x"ff"),
  1148 => (x"bf",x"97",x"d6",x"e3"),
  1149 => (x"74",x"87",x"d8",x"02"),
  1150 => (x"c1",x"91",x"de",x"49"),
  1151 => (x"e4",x"e8",x"c2",x"84"),
  1152 => (x"c2",x"83",x"71",x"4b"),
  1153 => (x"dd",x"4a",x"d6",x"e3"),
  1154 => (x"da",x"fa",x"fe",x"49"),
  1155 => (x"74",x"87",x"d8",x"87"),
  1156 => (x"c2",x"93",x"de",x"4b"),
  1157 => (x"cb",x"83",x"e4",x"e8"),
  1158 => (x"51",x"c0",x"49",x"a3"),
  1159 => (x"6e",x"73",x"84",x"c1"),
  1160 => (x"fe",x"49",x"cb",x"4a"),
  1161 => (x"c4",x"87",x"c0",x"fa"),
  1162 => (x"80",x"c1",x"48",x"66"),
  1163 => (x"c7",x"58",x"a6",x"c8"),
  1164 => (x"c5",x"c0",x"03",x"ac"),
  1165 => (x"fc",x"05",x"6e",x"87"),
  1166 => (x"48",x"74",x"87",x"e4"),
  1167 => (x"f6",x"f4",x"8e",x"f4"),
  1168 => (x"1e",x"73",x"1e",x"87"),
  1169 => (x"cb",x"49",x"4b",x"71"),
  1170 => (x"ec",x"e3",x"c1",x"91"),
  1171 => (x"4a",x"a1",x"c8",x"81"),
  1172 => (x"48",x"d8",x"e3",x"c1"),
  1173 => (x"a1",x"c9",x"50",x"12"),
  1174 => (x"ea",x"f8",x"c0",x"4a"),
  1175 => (x"ca",x"50",x"12",x"48"),
  1176 => (x"d9",x"e3",x"c1",x"81"),
  1177 => (x"c1",x"50",x"11",x"48"),
  1178 => (x"bf",x"97",x"d9",x"e3"),
  1179 => (x"49",x"c0",x"1e",x"49"),
  1180 => (x"c2",x"87",x"cb",x"f5"),
  1181 => (x"de",x"48",x"f8",x"e7"),
  1182 => (x"d6",x"49",x"c1",x"78"),
  1183 => (x"f3",x"26",x"87",x"c1"),
  1184 => (x"5e",x"0e",x"87",x"f9"),
  1185 => (x"0e",x"5d",x"5c",x"5b"),
  1186 => (x"4d",x"71",x"86",x"f4"),
  1187 => (x"c1",x"91",x"cb",x"49"),
  1188 => (x"c8",x"81",x"ec",x"e3"),
  1189 => (x"a1",x"ca",x"4a",x"a1"),
  1190 => (x"48",x"a6",x"c4",x"7e"),
  1191 => (x"bf",x"c0",x"ec",x"c2"),
  1192 => (x"bf",x"97",x"6e",x"78"),
  1193 => (x"48",x"66",x"c4",x"4b"),
  1194 => (x"4b",x"70",x"28",x"73"),
  1195 => (x"cc",x"48",x"12",x"4c"),
  1196 => (x"9c",x"70",x"58",x"a6"),
  1197 => (x"81",x"c9",x"84",x"c1"),
  1198 => (x"b7",x"49",x"69",x"97"),
  1199 => (x"87",x"c2",x"04",x"ac"),
  1200 => (x"97",x"6e",x"4c",x"c0"),
  1201 => (x"66",x"c8",x"4a",x"bf"),
  1202 => (x"ff",x"31",x"72",x"49"),
  1203 => (x"99",x"66",x"c4",x"b9"),
  1204 => (x"30",x"72",x"48",x"74"),
  1205 => (x"71",x"48",x"4a",x"70"),
  1206 => (x"c4",x"ec",x"c2",x"b0"),
  1207 => (x"f8",x"e4",x"c0",x"58"),
  1208 => (x"d4",x"49",x"c0",x"87"),
  1209 => (x"49",x"75",x"87",x"d9"),
  1210 => (x"87",x"ed",x"f6",x"c0"),
  1211 => (x"c6",x"f2",x"8e",x"f4"),
  1212 => (x"1e",x"73",x"1e",x"87"),
  1213 => (x"fe",x"49",x"4b",x"71"),
  1214 => (x"49",x"73",x"87",x"c8"),
  1215 => (x"f1",x"87",x"c3",x"fe"),
  1216 => (x"73",x"1e",x"87",x"f9"),
  1217 => (x"c6",x"4b",x"71",x"1e"),
  1218 => (x"c0",x"02",x"4a",x"a3"),
  1219 => (x"8a",x"c1",x"87",x"e3"),
  1220 => (x"8a",x"87",x"d6",x"02"),
  1221 => (x"87",x"e8",x"c1",x"02"),
  1222 => (x"ca",x"c1",x"02",x"8a"),
  1223 => (x"c0",x"02",x"8a",x"87"),
  1224 => (x"02",x"8a",x"87",x"ef"),
  1225 => (x"e9",x"c1",x"87",x"d9"),
  1226 => (x"f6",x"49",x"c7",x"87"),
  1227 => (x"ec",x"c1",x"87",x"c3"),
  1228 => (x"f8",x"e7",x"c2",x"87"),
  1229 => (x"c1",x"78",x"df",x"48"),
  1230 => (x"87",x"c3",x"d3",x"49"),
  1231 => (x"c2",x"87",x"de",x"c1"),
  1232 => (x"02",x"bf",x"d0",x"e8"),
  1233 => (x"48",x"87",x"cb",x"c1"),
  1234 => (x"e8",x"c2",x"88",x"c1"),
  1235 => (x"c1",x"c1",x"58",x"d4"),
  1236 => (x"d4",x"e8",x"c2",x"87"),
  1237 => (x"f9",x"c0",x"02",x"bf"),
  1238 => (x"d0",x"e8",x"c2",x"87"),
  1239 => (x"80",x"c1",x"48",x"bf"),
  1240 => (x"58",x"d4",x"e8",x"c2"),
  1241 => (x"c2",x"87",x"eb",x"c0"),
  1242 => (x"49",x"bf",x"d0",x"e8"),
  1243 => (x"e8",x"c2",x"89",x"c6"),
  1244 => (x"b7",x"c0",x"59",x"d4"),
  1245 => (x"87",x"da",x"03",x"a9"),
  1246 => (x"48",x"d0",x"e8",x"c2"),
  1247 => (x"87",x"d2",x"78",x"c0"),
  1248 => (x"bf",x"d4",x"e8",x"c2"),
  1249 => (x"c2",x"87",x"cb",x"02"),
  1250 => (x"48",x"bf",x"d0",x"e8"),
  1251 => (x"e8",x"c2",x"80",x"c6"),
  1252 => (x"49",x"c0",x"58",x"d4"),
  1253 => (x"73",x"87",x"e8",x"d1"),
  1254 => (x"fc",x"f3",x"c0",x"49"),
  1255 => (x"87",x"db",x"ef",x"87"),
  1256 => (x"5c",x"5b",x"5e",x"0e"),
  1257 => (x"d4",x"ff",x"0e",x"5d"),
  1258 => (x"59",x"a6",x"dc",x"86"),
  1259 => (x"c0",x"48",x"a6",x"c8"),
  1260 => (x"c1",x"80",x"c4",x"78"),
  1261 => (x"c4",x"78",x"66",x"c0"),
  1262 => (x"c4",x"78",x"c1",x"80"),
  1263 => (x"c2",x"78",x"c1",x"80"),
  1264 => (x"c1",x"48",x"d4",x"e8"),
  1265 => (x"f8",x"e7",x"c2",x"78"),
  1266 => (x"a8",x"de",x"48",x"bf"),
  1267 => (x"f4",x"87",x"c9",x"05"),
  1268 => (x"a6",x"cc",x"87",x"e6"),
  1269 => (x"87",x"e6",x"cf",x"58"),
  1270 => (x"e4",x"87",x"df",x"e3"),
  1271 => (x"ce",x"e3",x"87",x"c1"),
  1272 => (x"c0",x"4c",x"70",x"87"),
  1273 => (x"c1",x"02",x"ac",x"fb"),
  1274 => (x"66",x"d8",x"87",x"fb"),
  1275 => (x"87",x"ed",x"c1",x"05"),
  1276 => (x"4a",x"66",x"fc",x"c0"),
  1277 => (x"7e",x"6a",x"82",x"c4"),
  1278 => (x"df",x"c1",x"1e",x"72"),
  1279 => (x"66",x"c4",x"48",x"f3"),
  1280 => (x"4a",x"a1",x"c8",x"49"),
  1281 => (x"aa",x"71",x"41",x"20"),
  1282 => (x"10",x"87",x"f9",x"05"),
  1283 => (x"c0",x"4a",x"26",x"51"),
  1284 => (x"c1",x"48",x"66",x"fc"),
  1285 => (x"6a",x"78",x"c1",x"c9"),
  1286 => (x"74",x"81",x"c7",x"49"),
  1287 => (x"66",x"fc",x"c0",x"51"),
  1288 => (x"c1",x"81",x"c8",x"49"),
  1289 => (x"66",x"fc",x"c0",x"51"),
  1290 => (x"c0",x"81",x"c9",x"49"),
  1291 => (x"66",x"fc",x"c0",x"51"),
  1292 => (x"c0",x"81",x"ca",x"49"),
  1293 => (x"d8",x"1e",x"c1",x"51"),
  1294 => (x"c8",x"49",x"6a",x"1e"),
  1295 => (x"87",x"f3",x"e2",x"81"),
  1296 => (x"c0",x"c1",x"86",x"c8"),
  1297 => (x"a8",x"c0",x"48",x"66"),
  1298 => (x"c8",x"87",x"c7",x"01"),
  1299 => (x"78",x"c1",x"48",x"a6"),
  1300 => (x"c0",x"c1",x"87",x"ce"),
  1301 => (x"88",x"c1",x"48",x"66"),
  1302 => (x"c3",x"58",x"a6",x"d0"),
  1303 => (x"87",x"ff",x"e1",x"87"),
  1304 => (x"c2",x"48",x"a6",x"d0"),
  1305 => (x"02",x"9c",x"74",x"78"),
  1306 => (x"c8",x"87",x"cf",x"cd"),
  1307 => (x"c4",x"c1",x"48",x"66"),
  1308 => (x"cd",x"03",x"a8",x"66"),
  1309 => (x"a6",x"dc",x"87",x"c4"),
  1310 => (x"e8",x"78",x"c0",x"48"),
  1311 => (x"e0",x"78",x"c0",x"80"),
  1312 => (x"4c",x"70",x"87",x"ed"),
  1313 => (x"05",x"ac",x"d0",x"c1"),
  1314 => (x"c4",x"87",x"d7",x"c2"),
  1315 => (x"d1",x"e3",x"7e",x"66"),
  1316 => (x"58",x"a6",x"c8",x"87"),
  1317 => (x"70",x"87",x"d8",x"e0"),
  1318 => (x"ac",x"ec",x"c0",x"4c"),
  1319 => (x"87",x"ed",x"c1",x"05"),
  1320 => (x"cb",x"49",x"66",x"c8"),
  1321 => (x"66",x"fc",x"c0",x"91"),
  1322 => (x"4a",x"a1",x"c4",x"81"),
  1323 => (x"a1",x"c8",x"4d",x"6a"),
  1324 => (x"52",x"66",x"c4",x"4a"),
  1325 => (x"79",x"f1",x"c2",x"c1"),
  1326 => (x"87",x"f3",x"df",x"ff"),
  1327 => (x"02",x"9c",x"4c",x"70"),
  1328 => (x"fb",x"c0",x"87",x"d9"),
  1329 => (x"87",x"d3",x"02",x"ac"),
  1330 => (x"df",x"ff",x"55",x"74"),
  1331 => (x"4c",x"70",x"87",x"e1"),
  1332 => (x"87",x"c7",x"02",x"9c"),
  1333 => (x"05",x"ac",x"fb",x"c0"),
  1334 => (x"c0",x"87",x"ed",x"ff"),
  1335 => (x"c1",x"c2",x"55",x"e0"),
  1336 => (x"7d",x"97",x"c0",x"55"),
  1337 => (x"6e",x"48",x"66",x"d8"),
  1338 => (x"87",x"db",x"05",x"a8"),
  1339 => (x"cc",x"48",x"66",x"c8"),
  1340 => (x"ca",x"04",x"a8",x"66"),
  1341 => (x"48",x"66",x"c8",x"87"),
  1342 => (x"a6",x"cc",x"80",x"c1"),
  1343 => (x"cc",x"87",x"c8",x"58"),
  1344 => (x"88",x"c1",x"48",x"66"),
  1345 => (x"ff",x"58",x"a6",x"d0"),
  1346 => (x"70",x"87",x"e4",x"de"),
  1347 => (x"ac",x"d0",x"c1",x"4c"),
  1348 => (x"d4",x"87",x"c8",x"05"),
  1349 => (x"80",x"c1",x"48",x"66"),
  1350 => (x"c1",x"58",x"a6",x"d8"),
  1351 => (x"fd",x"02",x"ac",x"d0"),
  1352 => (x"66",x"c4",x"87",x"e9"),
  1353 => (x"a8",x"66",x"d8",x"48"),
  1354 => (x"87",x"e0",x"c9",x"05"),
  1355 => (x"48",x"a6",x"e0",x"c0"),
  1356 => (x"48",x"74",x"78",x"c0"),
  1357 => (x"70",x"88",x"fb",x"c0"),
  1358 => (x"02",x"98",x"48",x"7e"),
  1359 => (x"48",x"87",x"e2",x"c9"),
  1360 => (x"7e",x"70",x"88",x"cb"),
  1361 => (x"c1",x"02",x"98",x"48"),
  1362 => (x"c9",x"48",x"87",x"cd"),
  1363 => (x"48",x"7e",x"70",x"88"),
  1364 => (x"fe",x"c3",x"02",x"98"),
  1365 => (x"88",x"c4",x"48",x"87"),
  1366 => (x"98",x"48",x"7e",x"70"),
  1367 => (x"48",x"87",x"ce",x"02"),
  1368 => (x"7e",x"70",x"88",x"c1"),
  1369 => (x"c3",x"02",x"98",x"48"),
  1370 => (x"d6",x"c8",x"87",x"e9"),
  1371 => (x"48",x"a6",x"dc",x"87"),
  1372 => (x"ff",x"78",x"f0",x"c0"),
  1373 => (x"70",x"87",x"f8",x"dc"),
  1374 => (x"ac",x"ec",x"c0",x"4c"),
  1375 => (x"87",x"c4",x"c0",x"02"),
  1376 => (x"5c",x"a6",x"e0",x"c0"),
  1377 => (x"02",x"ac",x"ec",x"c0"),
  1378 => (x"dc",x"ff",x"87",x"cd"),
  1379 => (x"4c",x"70",x"87",x"e1"),
  1380 => (x"05",x"ac",x"ec",x"c0"),
  1381 => (x"c0",x"87",x"f3",x"ff"),
  1382 => (x"c0",x"02",x"ac",x"ec"),
  1383 => (x"dc",x"ff",x"87",x"c4"),
  1384 => (x"1e",x"c0",x"87",x"cd"),
  1385 => (x"66",x"d0",x"1e",x"ca"),
  1386 => (x"c1",x"91",x"cb",x"49"),
  1387 => (x"71",x"48",x"66",x"c4"),
  1388 => (x"58",x"a6",x"cc",x"80"),
  1389 => (x"c4",x"48",x"66",x"c8"),
  1390 => (x"58",x"a6",x"d0",x"80"),
  1391 => (x"49",x"bf",x"66",x"cc"),
  1392 => (x"87",x"ef",x"dc",x"ff"),
  1393 => (x"1e",x"de",x"1e",x"c1"),
  1394 => (x"49",x"bf",x"66",x"d4"),
  1395 => (x"87",x"e3",x"dc",x"ff"),
  1396 => (x"49",x"70",x"86",x"d0"),
  1397 => (x"88",x"08",x"c0",x"48"),
  1398 => (x"58",x"a6",x"e8",x"c0"),
  1399 => (x"c0",x"06",x"a8",x"c0"),
  1400 => (x"e4",x"c0",x"87",x"ee"),
  1401 => (x"a8",x"dd",x"48",x"66"),
  1402 => (x"87",x"e4",x"c0",x"03"),
  1403 => (x"49",x"bf",x"66",x"c4"),
  1404 => (x"81",x"66",x"e4",x"c0"),
  1405 => (x"c0",x"51",x"e0",x"c0"),
  1406 => (x"c1",x"49",x"66",x"e4"),
  1407 => (x"bf",x"66",x"c4",x"81"),
  1408 => (x"51",x"c1",x"c2",x"81"),
  1409 => (x"49",x"66",x"e4",x"c0"),
  1410 => (x"66",x"c4",x"81",x"c2"),
  1411 => (x"51",x"c0",x"81",x"bf"),
  1412 => (x"c9",x"c1",x"48",x"6e"),
  1413 => (x"49",x"6e",x"78",x"c1"),
  1414 => (x"66",x"d0",x"81",x"c8"),
  1415 => (x"c9",x"49",x"6e",x"51"),
  1416 => (x"51",x"66",x"d4",x"81"),
  1417 => (x"81",x"ca",x"49",x"6e"),
  1418 => (x"d0",x"51",x"66",x"dc"),
  1419 => (x"80",x"c1",x"48",x"66"),
  1420 => (x"c8",x"58",x"a6",x"d4"),
  1421 => (x"66",x"cc",x"48",x"66"),
  1422 => (x"cb",x"c0",x"04",x"a8"),
  1423 => (x"48",x"66",x"c8",x"87"),
  1424 => (x"a6",x"cc",x"80",x"c1"),
  1425 => (x"87",x"d9",x"c5",x"58"),
  1426 => (x"c1",x"48",x"66",x"cc"),
  1427 => (x"58",x"a6",x"d0",x"88"),
  1428 => (x"ff",x"87",x"ce",x"c5"),
  1429 => (x"c0",x"87",x"cb",x"dc"),
  1430 => (x"ff",x"58",x"a6",x"e8"),
  1431 => (x"c0",x"87",x"c3",x"dc"),
  1432 => (x"c0",x"58",x"a6",x"e0"),
  1433 => (x"c0",x"05",x"a8",x"ec"),
  1434 => (x"a6",x"dc",x"87",x"ca"),
  1435 => (x"66",x"e4",x"c0",x"48"),
  1436 => (x"87",x"c4",x"c0",x"78"),
  1437 => (x"87",x"f7",x"d8",x"ff"),
  1438 => (x"cb",x"49",x"66",x"c8"),
  1439 => (x"66",x"fc",x"c0",x"91"),
  1440 => (x"70",x"80",x"71",x"48"),
  1441 => (x"82",x"c8",x"4a",x"7e"),
  1442 => (x"81",x"ca",x"49",x"6e"),
  1443 => (x"51",x"66",x"e4",x"c0"),
  1444 => (x"c1",x"49",x"66",x"dc"),
  1445 => (x"66",x"e4",x"c0",x"81"),
  1446 => (x"71",x"48",x"c1",x"89"),
  1447 => (x"c1",x"49",x"70",x"30"),
  1448 => (x"7a",x"97",x"71",x"89"),
  1449 => (x"bf",x"c0",x"ec",x"c2"),
  1450 => (x"66",x"e4",x"c0",x"49"),
  1451 => (x"4a",x"6a",x"97",x"29"),
  1452 => (x"c0",x"98",x"71",x"48"),
  1453 => (x"6e",x"58",x"a6",x"ec"),
  1454 => (x"69",x"81",x"c4",x"49"),
  1455 => (x"48",x"66",x"d8",x"4d"),
  1456 => (x"02",x"a8",x"66",x"c4"),
  1457 => (x"c4",x"87",x"c8",x"c0"),
  1458 => (x"78",x"c0",x"48",x"a6"),
  1459 => (x"c4",x"87",x"c5",x"c0"),
  1460 => (x"78",x"c1",x"48",x"a6"),
  1461 => (x"c0",x"1e",x"66",x"c4"),
  1462 => (x"49",x"75",x"1e",x"e0"),
  1463 => (x"87",x"d3",x"d8",x"ff"),
  1464 => (x"4c",x"70",x"86",x"c8"),
  1465 => (x"06",x"ac",x"b7",x"c0"),
  1466 => (x"74",x"87",x"d4",x"c1"),
  1467 => (x"49",x"e0",x"c0",x"85"),
  1468 => (x"4b",x"75",x"89",x"74"),
  1469 => (x"4a",x"fc",x"df",x"c1"),
  1470 => (x"ea",x"e6",x"fe",x"71"),
  1471 => (x"c0",x"85",x"c2",x"87"),
  1472 => (x"c1",x"48",x"66",x"e0"),
  1473 => (x"a6",x"e4",x"c0",x"80"),
  1474 => (x"66",x"e8",x"c0",x"58"),
  1475 => (x"70",x"81",x"c1",x"49"),
  1476 => (x"c8",x"c0",x"02",x"a9"),
  1477 => (x"48",x"a6",x"c4",x"87"),
  1478 => (x"c5",x"c0",x"78",x"c0"),
  1479 => (x"48",x"a6",x"c4",x"87"),
  1480 => (x"66",x"c4",x"78",x"c1"),
  1481 => (x"49",x"a4",x"c2",x"1e"),
  1482 => (x"71",x"48",x"e0",x"c0"),
  1483 => (x"1e",x"49",x"70",x"88"),
  1484 => (x"d6",x"ff",x"49",x"75"),
  1485 => (x"86",x"c8",x"87",x"fd"),
  1486 => (x"01",x"a8",x"b7",x"c0"),
  1487 => (x"c0",x"87",x"c0",x"ff"),
  1488 => (x"c0",x"02",x"66",x"e0"),
  1489 => (x"49",x"6e",x"87",x"d1"),
  1490 => (x"e0",x"c0",x"81",x"c9"),
  1491 => (x"48",x"6e",x"51",x"66"),
  1492 => (x"78",x"c2",x"ca",x"c1"),
  1493 => (x"6e",x"87",x"cc",x"c0"),
  1494 => (x"c2",x"81",x"c9",x"49"),
  1495 => (x"c1",x"48",x"6e",x"51"),
  1496 => (x"c8",x"78",x"f1",x"cb"),
  1497 => (x"66",x"cc",x"48",x"66"),
  1498 => (x"cb",x"c0",x"04",x"a8"),
  1499 => (x"48",x"66",x"c8",x"87"),
  1500 => (x"a6",x"cc",x"80",x"c1"),
  1501 => (x"87",x"e9",x"c0",x"58"),
  1502 => (x"c1",x"48",x"66",x"cc"),
  1503 => (x"58",x"a6",x"d0",x"88"),
  1504 => (x"ff",x"87",x"de",x"c0"),
  1505 => (x"70",x"87",x"d8",x"d5"),
  1506 => (x"87",x"d5",x"c0",x"4c"),
  1507 => (x"05",x"ac",x"c6",x"c1"),
  1508 => (x"d0",x"87",x"c8",x"c0"),
  1509 => (x"80",x"c1",x"48",x"66"),
  1510 => (x"ff",x"58",x"a6",x"d4"),
  1511 => (x"70",x"87",x"c0",x"d5"),
  1512 => (x"48",x"66",x"d4",x"4c"),
  1513 => (x"a6",x"d8",x"80",x"c1"),
  1514 => (x"02",x"9c",x"74",x"58"),
  1515 => (x"c8",x"87",x"cb",x"c0"),
  1516 => (x"c4",x"c1",x"48",x"66"),
  1517 => (x"f2",x"04",x"a8",x"66"),
  1518 => (x"d4",x"ff",x"87",x"fc"),
  1519 => (x"66",x"c8",x"87",x"d8"),
  1520 => (x"03",x"a8",x"c7",x"48"),
  1521 => (x"c2",x"87",x"e5",x"c0"),
  1522 => (x"c0",x"48",x"d4",x"e8"),
  1523 => (x"49",x"66",x"c8",x"78"),
  1524 => (x"fc",x"c0",x"91",x"cb"),
  1525 => (x"a1",x"c4",x"81",x"66"),
  1526 => (x"c0",x"4a",x"6a",x"4a"),
  1527 => (x"66",x"c8",x"79",x"52"),
  1528 => (x"cc",x"80",x"c1",x"48"),
  1529 => (x"a8",x"c7",x"58",x"a6"),
  1530 => (x"87",x"db",x"ff",x"04"),
  1531 => (x"ff",x"8e",x"d4",x"ff"),
  1532 => (x"4c",x"87",x"c4",x"de"),
  1533 => (x"20",x"64",x"61",x"6f"),
  1534 => (x"00",x"20",x"2e",x"2a"),
  1535 => (x"1e",x"00",x"20",x"3a"),
  1536 => (x"4b",x"71",x"1e",x"73"),
  1537 => (x"87",x"c6",x"02",x"9b"),
  1538 => (x"48",x"d0",x"e8",x"c2"),
  1539 => (x"1e",x"c7",x"78",x"c0"),
  1540 => (x"bf",x"d0",x"e8",x"c2"),
  1541 => (x"ec",x"e3",x"c1",x"1e"),
  1542 => (x"f8",x"e7",x"c2",x"1e"),
  1543 => (x"ff",x"ed",x"49",x"bf"),
  1544 => (x"c2",x"86",x"cc",x"87"),
  1545 => (x"49",x"bf",x"f8",x"e7"),
  1546 => (x"73",x"87",x"e5",x"e2"),
  1547 => (x"87",x"c8",x"02",x"9b"),
  1548 => (x"49",x"ec",x"e3",x"c1"),
  1549 => (x"87",x"f3",x"e2",x"c0"),
  1550 => (x"87",x"ff",x"dc",x"ff"),
  1551 => (x"d8",x"e3",x"c1",x"1e"),
  1552 => (x"c1",x"50",x"c0",x"48"),
  1553 => (x"49",x"bf",x"cf",x"e5"),
  1554 => (x"87",x"df",x"d7",x"ff"),
  1555 => (x"4f",x"26",x"48",x"c0"),
  1556 => (x"87",x"df",x"c7",x"1e"),
  1557 => (x"e6",x"fe",x"49",x"c1"),
  1558 => (x"f6",x"e9",x"fe",x"87"),
  1559 => (x"02",x"98",x"70",x"87"),
  1560 => (x"f2",x"fe",x"87",x"cd"),
  1561 => (x"98",x"70",x"87",x"f0"),
  1562 => (x"c1",x"87",x"c4",x"02"),
  1563 => (x"c0",x"87",x"c2",x"4a"),
  1564 => (x"05",x"9a",x"72",x"4a"),
  1565 => (x"1e",x"c0",x"87",x"ce"),
  1566 => (x"49",x"eb",x"e2",x"c1"),
  1567 => (x"87",x"de",x"ef",x"c0"),
  1568 => (x"87",x"fe",x"86",x"c4"),
  1569 => (x"48",x"d0",x"e8",x"c2"),
  1570 => (x"e7",x"c2",x"78",x"c0"),
  1571 => (x"78",x"c0",x"48",x"f8"),
  1572 => (x"f6",x"e2",x"c1",x"1e"),
  1573 => (x"c5",x"ef",x"c0",x"49"),
  1574 => (x"fe",x"1e",x"c0",x"87"),
  1575 => (x"49",x"70",x"87",x"de"),
  1576 => (x"87",x"fa",x"ee",x"c0"),
  1577 => (x"f8",x"87",x"cb",x"c3"),
  1578 => (x"53",x"4f",x"26",x"8e"),
  1579 => (x"61",x"66",x"20",x"44"),
  1580 => (x"64",x"65",x"6c",x"69"),
  1581 => (x"6f",x"42",x"00",x"2e"),
  1582 => (x"6e",x"69",x"74",x"6f"),
  1583 => (x"2e",x"2e",x"2e",x"67"),
  1584 => (x"e2",x"c0",x"1e",x"00"),
  1585 => (x"f2",x"c0",x"87",x"e2"),
  1586 => (x"87",x"f6",x"87",x"ce"),
  1587 => (x"fd",x"1e",x"4f",x"26"),
  1588 => (x"87",x"ed",x"87",x"fe"),
  1589 => (x"4f",x"26",x"48",x"c0"),
  1590 => (x"00",x"01",x"00",x"00"),
  1591 => (x"20",x"80",x"00",x"00"),
  1592 => (x"74",x"69",x"78",x"45"),
  1593 => (x"42",x"20",x"80",x"00"),
  1594 => (x"00",x"6b",x"63",x"61"),
  1595 => (x"00",x"00",x"0f",x"fe"),
  1596 => (x"00",x"00",x"2a",x"24"),
  1597 => (x"fe",x"00",x"00",x"00"),
  1598 => (x"42",x"00",x"00",x"0f"),
  1599 => (x"00",x"00",x"00",x"2a"),
  1600 => (x"0f",x"fe",x"00",x"00"),
  1601 => (x"2a",x"60",x"00",x"00"),
  1602 => (x"00",x"00",x"00",x"00"),
  1603 => (x"00",x"0f",x"fe",x"00"),
  1604 => (x"00",x"2a",x"7e",x"00"),
  1605 => (x"00",x"00",x"00",x"00"),
  1606 => (x"00",x"00",x"0f",x"fe"),
  1607 => (x"00",x"00",x"2a",x"9c"),
  1608 => (x"fe",x"00",x"00",x"00"),
  1609 => (x"ba",x"00",x"00",x"0f"),
  1610 => (x"00",x"00",x"00",x"2a"),
  1611 => (x"0f",x"fe",x"00",x"00"),
  1612 => (x"2a",x"d8",x"00",x"00"),
  1613 => (x"00",x"00",x"00",x"00"),
  1614 => (x"00",x"10",x"b1",x"00"),
  1615 => (x"00",x"00",x"00",x"00"),
  1616 => (x"00",x"00",x"00",x"00"),
  1617 => (x"00",x"00",x"13",x"02"),
  1618 => (x"00",x"00",x"00",x"00"),
  1619 => (x"53",x"00",x"00",x"00"),
  1620 => (x"42",x"00",x"00",x"19"),
  1621 => (x"20",x"54",x"4f",x"4f"),
  1622 => (x"52",x"20",x"20",x"20"),
  1623 => (x"1e",x"00",x"4d",x"4f"),
  1624 => (x"c0",x"48",x"f0",x"fe"),
  1625 => (x"79",x"09",x"cd",x"78"),
  1626 => (x"1e",x"4f",x"26",x"09"),
  1627 => (x"48",x"bf",x"f0",x"fe"),
  1628 => (x"fe",x"1e",x"4f",x"26"),
  1629 => (x"78",x"c1",x"48",x"f0"),
  1630 => (x"fe",x"1e",x"4f",x"26"),
  1631 => (x"78",x"c0",x"48",x"f0"),
  1632 => (x"71",x"1e",x"4f",x"26"),
  1633 => (x"51",x"52",x"c0",x"4a"),
  1634 => (x"5e",x"0e",x"4f",x"26"),
  1635 => (x"0e",x"5d",x"5c",x"5b"),
  1636 => (x"4d",x"71",x"86",x"f4"),
  1637 => (x"c1",x"7e",x"6d",x"97"),
  1638 => (x"6c",x"97",x"4c",x"a5"),
  1639 => (x"58",x"a6",x"c8",x"48"),
  1640 => (x"66",x"c4",x"48",x"6e"),
  1641 => (x"87",x"c5",x"05",x"a8"),
  1642 => (x"e6",x"c0",x"48",x"ff"),
  1643 => (x"87",x"ca",x"ff",x"87"),
  1644 => (x"97",x"49",x"a5",x"c2"),
  1645 => (x"a3",x"71",x"4b",x"6c"),
  1646 => (x"4b",x"6b",x"97",x"4b"),
  1647 => (x"6e",x"7e",x"6c",x"97"),
  1648 => (x"c8",x"80",x"c1",x"48"),
  1649 => (x"98",x"c7",x"58",x"a6"),
  1650 => (x"70",x"58",x"a6",x"cc"),
  1651 => (x"e1",x"fe",x"7c",x"97"),
  1652 => (x"f4",x"48",x"73",x"87"),
  1653 => (x"26",x"4d",x"26",x"8e"),
  1654 => (x"26",x"4b",x"26",x"4c"),
  1655 => (x"5b",x"5e",x"0e",x"4f"),
  1656 => (x"86",x"f4",x"0e",x"5c"),
  1657 => (x"66",x"d8",x"4c",x"71"),
  1658 => (x"9a",x"ff",x"c3",x"4a"),
  1659 => (x"97",x"4b",x"a4",x"c2"),
  1660 => (x"a1",x"73",x"49",x"6c"),
  1661 => (x"97",x"51",x"72",x"49"),
  1662 => (x"48",x"6e",x"7e",x"6c"),
  1663 => (x"a6",x"c8",x"80",x"c1"),
  1664 => (x"cc",x"98",x"c7",x"58"),
  1665 => (x"54",x"70",x"58",x"a6"),
  1666 => (x"ca",x"ff",x"8e",x"f4"),
  1667 => (x"fd",x"1e",x"1e",x"87"),
  1668 => (x"bf",x"e0",x"87",x"e8"),
  1669 => (x"e0",x"c0",x"49",x"4a"),
  1670 => (x"cb",x"02",x"99",x"c0"),
  1671 => (x"c2",x"1e",x"72",x"87"),
  1672 => (x"fe",x"49",x"f6",x"eb"),
  1673 => (x"86",x"c4",x"87",x"f7"),
  1674 => (x"70",x"87",x"c0",x"fd"),
  1675 => (x"87",x"c2",x"fd",x"7e"),
  1676 => (x"1e",x"4f",x"26",x"26"),
  1677 => (x"49",x"f6",x"eb",x"c2"),
  1678 => (x"c1",x"87",x"c7",x"fd"),
  1679 => (x"fc",x"49",x"cd",x"e8"),
  1680 => (x"ee",x"c3",x"87",x"dd"),
  1681 => (x"0e",x"4f",x"26",x"87"),
  1682 => (x"5d",x"5c",x"5b",x"5e"),
  1683 => (x"c2",x"4d",x"71",x"0e"),
  1684 => (x"fc",x"49",x"f6",x"eb"),
  1685 => (x"4b",x"70",x"87",x"f4"),
  1686 => (x"04",x"ab",x"b7",x"c0"),
  1687 => (x"c3",x"87",x"c2",x"c3"),
  1688 => (x"c9",x"05",x"ab",x"f0"),
  1689 => (x"eb",x"ec",x"c1",x"87"),
  1690 => (x"c2",x"78",x"c1",x"48"),
  1691 => (x"e0",x"c3",x"87",x"e3"),
  1692 => (x"87",x"c9",x"05",x"ab"),
  1693 => (x"48",x"ef",x"ec",x"c1"),
  1694 => (x"d4",x"c2",x"78",x"c1"),
  1695 => (x"ef",x"ec",x"c1",x"87"),
  1696 => (x"87",x"c6",x"02",x"bf"),
  1697 => (x"4c",x"a3",x"c0",x"c2"),
  1698 => (x"4c",x"73",x"87",x"c2"),
  1699 => (x"bf",x"eb",x"ec",x"c1"),
  1700 => (x"87",x"e0",x"c0",x"02"),
  1701 => (x"b7",x"c4",x"49",x"74"),
  1702 => (x"ee",x"c1",x"91",x"29"),
  1703 => (x"4a",x"74",x"81",x"c2"),
  1704 => (x"92",x"c2",x"9a",x"cf"),
  1705 => (x"30",x"72",x"48",x"c1"),
  1706 => (x"ba",x"ff",x"4a",x"70"),
  1707 => (x"98",x"69",x"48",x"72"),
  1708 => (x"87",x"db",x"79",x"70"),
  1709 => (x"b7",x"c4",x"49",x"74"),
  1710 => (x"ee",x"c1",x"91",x"29"),
  1711 => (x"4a",x"74",x"81",x"c2"),
  1712 => (x"92",x"c2",x"9a",x"cf"),
  1713 => (x"30",x"72",x"48",x"c3"),
  1714 => (x"69",x"48",x"4a",x"70"),
  1715 => (x"75",x"79",x"70",x"b0"),
  1716 => (x"f0",x"c0",x"05",x"9d"),
  1717 => (x"48",x"d0",x"ff",x"87"),
  1718 => (x"ff",x"78",x"e1",x"c8"),
  1719 => (x"78",x"c5",x"48",x"d4"),
  1720 => (x"bf",x"ef",x"ec",x"c1"),
  1721 => (x"c3",x"87",x"c3",x"02"),
  1722 => (x"ec",x"c1",x"78",x"e0"),
  1723 => (x"c6",x"02",x"bf",x"eb"),
  1724 => (x"48",x"d4",x"ff",x"87"),
  1725 => (x"ff",x"78",x"f0",x"c3"),
  1726 => (x"0b",x"7b",x"0b",x"d4"),
  1727 => (x"c8",x"48",x"d0",x"ff"),
  1728 => (x"e0",x"c0",x"78",x"e1"),
  1729 => (x"ef",x"ec",x"c1",x"78"),
  1730 => (x"c1",x"78",x"c0",x"48"),
  1731 => (x"c0",x"48",x"eb",x"ec"),
  1732 => (x"f6",x"eb",x"c2",x"78"),
  1733 => (x"87",x"f2",x"f9",x"49"),
  1734 => (x"b7",x"c0",x"4b",x"70"),
  1735 => (x"fe",x"fc",x"03",x"ab"),
  1736 => (x"26",x"48",x"c0",x"87"),
  1737 => (x"26",x"4c",x"26",x"4d"),
  1738 => (x"00",x"4f",x"26",x"4b"),
  1739 => (x"00",x"00",x"00",x"00"),
  1740 => (x"1e",x"00",x"00",x"00"),
  1741 => (x"49",x"72",x"4a",x"c0"),
  1742 => (x"ee",x"c1",x"91",x"c4"),
  1743 => (x"79",x"c0",x"81",x"c2"),
  1744 => (x"b7",x"d0",x"82",x"c1"),
  1745 => (x"87",x"ee",x"04",x"aa"),
  1746 => (x"5e",x"0e",x"4f",x"26"),
  1747 => (x"0e",x"5d",x"5c",x"5b"),
  1748 => (x"e5",x"f8",x"4d",x"71"),
  1749 => (x"c4",x"4a",x"75",x"87"),
  1750 => (x"c1",x"92",x"2a",x"b7"),
  1751 => (x"75",x"82",x"c2",x"ee"),
  1752 => (x"c2",x"9c",x"cf",x"4c"),
  1753 => (x"4b",x"49",x"6a",x"94"),
  1754 => (x"9b",x"c3",x"2b",x"74"),
  1755 => (x"30",x"74",x"48",x"c2"),
  1756 => (x"bc",x"ff",x"4c",x"70"),
  1757 => (x"98",x"71",x"48",x"74"),
  1758 => (x"f5",x"f7",x"7a",x"70"),
  1759 => (x"fe",x"48",x"73",x"87"),
  1760 => (x"00",x"00",x"87",x"e1"),
  1761 => (x"00",x"00",x"00",x"00"),
  1762 => (x"00",x"00",x"00",x"00"),
  1763 => (x"00",x"00",x"00",x"00"),
  1764 => (x"00",x"00",x"00",x"00"),
  1765 => (x"00",x"00",x"00",x"00"),
  1766 => (x"00",x"00",x"00",x"00"),
  1767 => (x"00",x"00",x"00",x"00"),
  1768 => (x"00",x"00",x"00",x"00"),
  1769 => (x"00",x"00",x"00",x"00"),
  1770 => (x"00",x"00",x"00",x"00"),
  1771 => (x"00",x"00",x"00",x"00"),
  1772 => (x"00",x"00",x"00",x"00"),
  1773 => (x"00",x"00",x"00",x"00"),
  1774 => (x"00",x"00",x"00",x"00"),
  1775 => (x"00",x"00",x"00",x"00"),
  1776 => (x"ff",x"1e",x"00",x"00"),
  1777 => (x"e1",x"c8",x"48",x"d0"),
  1778 => (x"ff",x"48",x"71",x"78"),
  1779 => (x"26",x"78",x"08",x"d4"),
  1780 => (x"d0",x"ff",x"1e",x"4f"),
  1781 => (x"78",x"e1",x"c8",x"48"),
  1782 => (x"d4",x"ff",x"48",x"71"),
  1783 => (x"66",x"c4",x"78",x"08"),
  1784 => (x"08",x"d4",x"ff",x"48"),
  1785 => (x"1e",x"4f",x"26",x"78"),
  1786 => (x"66",x"c4",x"4a",x"71"),
  1787 => (x"49",x"72",x"1e",x"49"),
  1788 => (x"ff",x"87",x"de",x"ff"),
  1789 => (x"e0",x"c0",x"48",x"d0"),
  1790 => (x"4f",x"26",x"26",x"78"),
  1791 => (x"71",x"1e",x"73",x"1e"),
  1792 => (x"49",x"66",x"c8",x"4b"),
  1793 => (x"c1",x"4a",x"73",x"1e"),
  1794 => (x"ff",x"49",x"a2",x"e0"),
  1795 => (x"c4",x"26",x"87",x"d9"),
  1796 => (x"26",x"4d",x"26",x"87"),
  1797 => (x"26",x"4b",x"26",x"4c"),
  1798 => (x"d4",x"ff",x"1e",x"4f"),
  1799 => (x"7a",x"ff",x"c3",x"4a"),
  1800 => (x"c0",x"48",x"d0",x"ff"),
  1801 => (x"7a",x"de",x"78",x"e1"),
  1802 => (x"bf",x"c0",x"ec",x"c2"),
  1803 => (x"c8",x"48",x"49",x"7a"),
  1804 => (x"71",x"7a",x"70",x"28"),
  1805 => (x"70",x"28",x"d0",x"48"),
  1806 => (x"d8",x"48",x"71",x"7a"),
  1807 => (x"ff",x"7a",x"70",x"28"),
  1808 => (x"e0",x"c0",x"48",x"d0"),
  1809 => (x"1e",x"4f",x"26",x"78"),
  1810 => (x"c8",x"48",x"d0",x"ff"),
  1811 => (x"48",x"71",x"78",x"c9"),
  1812 => (x"78",x"08",x"d4",x"ff"),
  1813 => (x"71",x"1e",x"4f",x"26"),
  1814 => (x"87",x"eb",x"49",x"4a"),
  1815 => (x"c8",x"48",x"d0",x"ff"),
  1816 => (x"1e",x"4f",x"26",x"78"),
  1817 => (x"4b",x"71",x"1e",x"73"),
  1818 => (x"bf",x"d0",x"ec",x"c2"),
  1819 => (x"c2",x"87",x"c3",x"02"),
  1820 => (x"d0",x"ff",x"87",x"eb"),
  1821 => (x"78",x"c9",x"c8",x"48"),
  1822 => (x"e0",x"c0",x"48",x"73"),
  1823 => (x"08",x"d4",x"ff",x"b0"),
  1824 => (x"c4",x"ec",x"c2",x"78"),
  1825 => (x"c8",x"78",x"c0",x"48"),
  1826 => (x"87",x"c5",x"02",x"66"),
  1827 => (x"c2",x"49",x"ff",x"c3"),
  1828 => (x"c2",x"49",x"c0",x"87"),
  1829 => (x"cc",x"59",x"cc",x"ec"),
  1830 => (x"87",x"c6",x"02",x"66"),
  1831 => (x"4a",x"d5",x"d5",x"c5"),
  1832 => (x"ff",x"cf",x"87",x"c4"),
  1833 => (x"ec",x"c2",x"4a",x"ff"),
  1834 => (x"ec",x"c2",x"5a",x"d0"),
  1835 => (x"78",x"c1",x"48",x"d0"),
  1836 => (x"4d",x"26",x"87",x"c4"),
  1837 => (x"4b",x"26",x"4c",x"26"),
  1838 => (x"5e",x"0e",x"4f",x"26"),
  1839 => (x"0e",x"5d",x"5c",x"5b"),
  1840 => (x"ec",x"c2",x"4a",x"71"),
  1841 => (x"72",x"4c",x"bf",x"cc"),
  1842 => (x"87",x"cb",x"02",x"9a"),
  1843 => (x"c1",x"91",x"c8",x"49"),
  1844 => (x"71",x"4b",x"d9",x"f1"),
  1845 => (x"c1",x"87",x"c4",x"83"),
  1846 => (x"c0",x"4b",x"d9",x"f5"),
  1847 => (x"74",x"49",x"13",x"4d"),
  1848 => (x"c8",x"ec",x"c2",x"99"),
  1849 => (x"b8",x"71",x"48",x"bf"),
  1850 => (x"78",x"08",x"d4",x"ff"),
  1851 => (x"85",x"2c",x"b7",x"c1"),
  1852 => (x"04",x"ad",x"b7",x"c8"),
  1853 => (x"ec",x"c2",x"87",x"e7"),
  1854 => (x"c8",x"48",x"bf",x"c4"),
  1855 => (x"c8",x"ec",x"c2",x"80"),
  1856 => (x"87",x"ee",x"fe",x"58"),
  1857 => (x"71",x"1e",x"73",x"1e"),
  1858 => (x"9a",x"4a",x"13",x"4b"),
  1859 => (x"72",x"87",x"cb",x"02"),
  1860 => (x"87",x"e6",x"fe",x"49"),
  1861 => (x"05",x"9a",x"4a",x"13"),
  1862 => (x"d9",x"fe",x"87",x"f5"),
  1863 => (x"ec",x"c2",x"1e",x"87"),
  1864 => (x"c2",x"49",x"bf",x"c4"),
  1865 => (x"c1",x"48",x"c4",x"ec"),
  1866 => (x"c0",x"c4",x"78",x"a1"),
  1867 => (x"db",x"03",x"a9",x"b7"),
  1868 => (x"48",x"d4",x"ff",x"87"),
  1869 => (x"bf",x"c8",x"ec",x"c2"),
  1870 => (x"c4",x"ec",x"c2",x"78"),
  1871 => (x"ec",x"c2",x"49",x"bf"),
  1872 => (x"a1",x"c1",x"48",x"c4"),
  1873 => (x"b7",x"c0",x"c4",x"78"),
  1874 => (x"87",x"e5",x"04",x"a9"),
  1875 => (x"c8",x"48",x"d0",x"ff"),
  1876 => (x"d0",x"ec",x"c2",x"78"),
  1877 => (x"26",x"78",x"c0",x"48"),
  1878 => (x"00",x"00",x"00",x"4f"),
  1879 => (x"00",x"00",x"00",x"00"),
  1880 => (x"00",x"00",x"00",x"00"),
  1881 => (x"00",x"00",x"5f",x"5f"),
  1882 => (x"03",x"03",x"00",x"00"),
  1883 => (x"00",x"03",x"03",x"00"),
  1884 => (x"7f",x"7f",x"14",x"00"),
  1885 => (x"14",x"7f",x"7f",x"14"),
  1886 => (x"2e",x"24",x"00",x"00"),
  1887 => (x"12",x"3a",x"6b",x"6b"),
  1888 => (x"36",x"6a",x"4c",x"00"),
  1889 => (x"32",x"56",x"6c",x"18"),
  1890 => (x"4f",x"7e",x"30",x"00"),
  1891 => (x"68",x"3a",x"77",x"59"),
  1892 => (x"04",x"00",x"00",x"40"),
  1893 => (x"00",x"00",x"03",x"07"),
  1894 => (x"1c",x"00",x"00",x"00"),
  1895 => (x"00",x"41",x"63",x"3e"),
  1896 => (x"41",x"00",x"00",x"00"),
  1897 => (x"00",x"1c",x"3e",x"63"),
  1898 => (x"3e",x"2a",x"08",x"00"),
  1899 => (x"2a",x"3e",x"1c",x"1c"),
  1900 => (x"08",x"08",x"00",x"08"),
  1901 => (x"08",x"08",x"3e",x"3e"),
  1902 => (x"80",x"00",x"00",x"00"),
  1903 => (x"00",x"00",x"60",x"e0"),
  1904 => (x"08",x"08",x"00",x"00"),
  1905 => (x"08",x"08",x"08",x"08"),
  1906 => (x"00",x"00",x"00",x"00"),
  1907 => (x"00",x"00",x"60",x"60"),
  1908 => (x"30",x"60",x"40",x"00"),
  1909 => (x"03",x"06",x"0c",x"18"),
  1910 => (x"7f",x"3e",x"00",x"01"),
  1911 => (x"3e",x"7f",x"4d",x"59"),
  1912 => (x"06",x"04",x"00",x"00"),
  1913 => (x"00",x"00",x"7f",x"7f"),
  1914 => (x"63",x"42",x"00",x"00"),
  1915 => (x"46",x"4f",x"59",x"71"),
  1916 => (x"63",x"22",x"00",x"00"),
  1917 => (x"36",x"7f",x"49",x"49"),
  1918 => (x"16",x"1c",x"18",x"00"),
  1919 => (x"10",x"7f",x"7f",x"13"),
  1920 => (x"67",x"27",x"00",x"00"),
  1921 => (x"39",x"7d",x"45",x"45"),
  1922 => (x"7e",x"3c",x"00",x"00"),
  1923 => (x"30",x"79",x"49",x"4b"),
  1924 => (x"01",x"01",x"00",x"00"),
  1925 => (x"07",x"0f",x"79",x"71"),
  1926 => (x"7f",x"36",x"00",x"00"),
  1927 => (x"36",x"7f",x"49",x"49"),
  1928 => (x"4f",x"06",x"00",x"00"),
  1929 => (x"1e",x"3f",x"69",x"49"),
  1930 => (x"00",x"00",x"00",x"00"),
  1931 => (x"00",x"00",x"66",x"66"),
  1932 => (x"80",x"00",x"00",x"00"),
  1933 => (x"00",x"00",x"66",x"e6"),
  1934 => (x"08",x"08",x"00",x"00"),
  1935 => (x"22",x"22",x"14",x"14"),
  1936 => (x"14",x"14",x"00",x"00"),
  1937 => (x"14",x"14",x"14",x"14"),
  1938 => (x"22",x"22",x"00",x"00"),
  1939 => (x"08",x"08",x"14",x"14"),
  1940 => (x"03",x"02",x"00",x"00"),
  1941 => (x"06",x"0f",x"59",x"51"),
  1942 => (x"41",x"7f",x"3e",x"00"),
  1943 => (x"1e",x"1f",x"55",x"5d"),
  1944 => (x"7f",x"7e",x"00",x"00"),
  1945 => (x"7e",x"7f",x"09",x"09"),
  1946 => (x"7f",x"7f",x"00",x"00"),
  1947 => (x"36",x"7f",x"49",x"49"),
  1948 => (x"3e",x"1c",x"00",x"00"),
  1949 => (x"41",x"41",x"41",x"63"),
  1950 => (x"7f",x"7f",x"00",x"00"),
  1951 => (x"1c",x"3e",x"63",x"41"),
  1952 => (x"7f",x"7f",x"00",x"00"),
  1953 => (x"41",x"41",x"49",x"49"),
  1954 => (x"7f",x"7f",x"00",x"00"),
  1955 => (x"01",x"01",x"09",x"09"),
  1956 => (x"7f",x"3e",x"00",x"00"),
  1957 => (x"7a",x"7b",x"49",x"41"),
  1958 => (x"7f",x"7f",x"00",x"00"),
  1959 => (x"7f",x"7f",x"08",x"08"),
  1960 => (x"41",x"00",x"00",x"00"),
  1961 => (x"00",x"41",x"7f",x"7f"),
  1962 => (x"60",x"20",x"00",x"00"),
  1963 => (x"3f",x"7f",x"40",x"40"),
  1964 => (x"08",x"7f",x"7f",x"00"),
  1965 => (x"41",x"63",x"36",x"1c"),
  1966 => (x"7f",x"7f",x"00",x"00"),
  1967 => (x"40",x"40",x"40",x"40"),
  1968 => (x"06",x"7f",x"7f",x"00"),
  1969 => (x"7f",x"7f",x"06",x"0c"),
  1970 => (x"06",x"7f",x"7f",x"00"),
  1971 => (x"7f",x"7f",x"18",x"0c"),
  1972 => (x"7f",x"3e",x"00",x"00"),
  1973 => (x"3e",x"7f",x"41",x"41"),
  1974 => (x"7f",x"7f",x"00",x"00"),
  1975 => (x"06",x"0f",x"09",x"09"),
  1976 => (x"41",x"7f",x"3e",x"00"),
  1977 => (x"40",x"7e",x"7f",x"61"),
  1978 => (x"7f",x"7f",x"00",x"00"),
  1979 => (x"66",x"7f",x"19",x"09"),
  1980 => (x"6f",x"26",x"00",x"00"),
  1981 => (x"32",x"7b",x"59",x"4d"),
  1982 => (x"01",x"01",x"00",x"00"),
  1983 => (x"01",x"01",x"7f",x"7f"),
  1984 => (x"7f",x"3f",x"00",x"00"),
  1985 => (x"3f",x"7f",x"40",x"40"),
  1986 => (x"3f",x"0f",x"00",x"00"),
  1987 => (x"0f",x"3f",x"70",x"70"),
  1988 => (x"30",x"7f",x"7f",x"00"),
  1989 => (x"7f",x"7f",x"30",x"18"),
  1990 => (x"36",x"63",x"41",x"00"),
  1991 => (x"63",x"36",x"1c",x"1c"),
  1992 => (x"06",x"03",x"01",x"41"),
  1993 => (x"03",x"06",x"7c",x"7c"),
  1994 => (x"59",x"71",x"61",x"01"),
  1995 => (x"41",x"43",x"47",x"4d"),
  1996 => (x"7f",x"00",x"00",x"00"),
  1997 => (x"00",x"41",x"41",x"7f"),
  1998 => (x"06",x"03",x"01",x"00"),
  1999 => (x"60",x"30",x"18",x"0c"),
  2000 => (x"41",x"00",x"00",x"40"),
  2001 => (x"00",x"7f",x"7f",x"41"),
  2002 => (x"06",x"0c",x"08",x"00"),
  2003 => (x"08",x"0c",x"06",x"03"),
  2004 => (x"80",x"80",x"80",x"00"),
  2005 => (x"80",x"80",x"80",x"80"),
  2006 => (x"00",x"00",x"00",x"00"),
  2007 => (x"00",x"04",x"07",x"03"),
  2008 => (x"74",x"20",x"00",x"00"),
  2009 => (x"78",x"7c",x"54",x"54"),
  2010 => (x"7f",x"7f",x"00",x"00"),
  2011 => (x"38",x"7c",x"44",x"44"),
  2012 => (x"7c",x"38",x"00",x"00"),
  2013 => (x"00",x"44",x"44",x"44"),
  2014 => (x"7c",x"38",x"00",x"00"),
  2015 => (x"7f",x"7f",x"44",x"44"),
  2016 => (x"7c",x"38",x"00",x"00"),
  2017 => (x"18",x"5c",x"54",x"54"),
  2018 => (x"7e",x"04",x"00",x"00"),
  2019 => (x"00",x"05",x"05",x"7f"),
  2020 => (x"bc",x"18",x"00",x"00"),
  2021 => (x"7c",x"fc",x"a4",x"a4"),
  2022 => (x"7f",x"7f",x"00",x"00"),
  2023 => (x"78",x"7c",x"04",x"04"),
  2024 => (x"00",x"00",x"00",x"00"),
  2025 => (x"00",x"40",x"7d",x"3d"),
  2026 => (x"80",x"80",x"00",x"00"),
  2027 => (x"00",x"7d",x"fd",x"80"),
  2028 => (x"7f",x"7f",x"00",x"00"),
  2029 => (x"44",x"6c",x"38",x"10"),
  2030 => (x"00",x"00",x"00",x"00"),
  2031 => (x"00",x"40",x"7f",x"3f"),
  2032 => (x"0c",x"7c",x"7c",x"00"),
  2033 => (x"78",x"7c",x"0c",x"18"),
  2034 => (x"7c",x"7c",x"00",x"00"),
  2035 => (x"78",x"7c",x"04",x"04"),
  2036 => (x"7c",x"38",x"00",x"00"),
  2037 => (x"38",x"7c",x"44",x"44"),
  2038 => (x"fc",x"fc",x"00",x"00"),
  2039 => (x"18",x"3c",x"24",x"24"),
  2040 => (x"3c",x"18",x"00",x"00"),
  2041 => (x"fc",x"fc",x"24",x"24"),
  2042 => (x"7c",x"7c",x"00",x"00"),
  2043 => (x"08",x"0c",x"04",x"04"),
  2044 => (x"5c",x"48",x"00",x"00"),
  2045 => (x"20",x"74",x"54",x"54"),
  2046 => (x"3f",x"04",x"00",x"00"),
  2047 => (x"00",x"44",x"44",x"7f"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

