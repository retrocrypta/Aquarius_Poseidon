library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom1 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom1 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"c8edc287",
    12 => x"86c0c84e",
    13 => x"49c8edc2",
    14 => x"48e0dac2",
    15 => x"4040c089",
    16 => x"89d04040",
    17 => x"c187f603",
    18 => x"0087c3e2",
    19 => x"721e87fd",
    20 => x"121e731e",
    21 => x"ca021148",
    22 => x"dfc34b87",
    23 => x"88739b98",
    24 => x"2687f002",
    25 => x"264a264b",
    26 => x"1e731e4f",
    27 => x"8bc11e72",
    28 => x"1287ca04",
    29 => x"c4021148",
    30 => x"f1028887",
    31 => x"264a2687",
    32 => x"1e4f264b",
    33 => x"1e731e74",
    34 => x"8bc11e72",
    35 => x"1287d004",
    36 => x"ca021148",
    37 => x"dfc34c87",
    38 => x"88749c98",
    39 => x"2687eb02",
    40 => x"264b264a",
    41 => x"1e4f264c",
    42 => x"73814873",
    43 => x"87c502a9",
    44 => x"f6055312",
    45 => x"1e4f2687",
    46 => x"66c44a71",
    47 => x"88c14849",
    48 => x"7158a6c8",
    49 => x"87d40299",
    50 => x"d4ff4812",
    51 => x"66c47808",
    52 => x"88c14849",
    53 => x"7158a6c8",
    54 => x"87ec0599",
    55 => x"711e4f26",
    56 => x"4966c44a",
    57 => x"c888c148",
    58 => x"997158a6",
    59 => x"ff87d602",
    60 => x"ffc348d4",
    61 => x"c4526878",
    62 => x"c1484966",
    63 => x"58a6c888",
    64 => x"ea059971",
    65 => x"1e4f2687",
    66 => x"d4ff1e73",
    67 => x"7bffc34b",
    68 => x"ffc34a6b",
    69 => x"c8496b7b",
    70 => x"c3b17232",
    71 => x"4a6b7bff",
    72 => x"b27131c8",
    73 => x"6b7bffc3",
    74 => x"7232c849",
    75 => x"c44871b1",
    76 => x"264d2687",
    77 => x"264b264c",
    78 => x"5b5e0e4f",
    79 => x"710e5d5c",
    80 => x"4cd4ff4a",
    81 => x"ffc34872",
    82 => x"c27c7098",
    83 => x"05bfe0da",
    84 => x"66d087c8",
    85 => x"d430c948",
    86 => x"66d058a6",
    87 => x"7129d849",
    88 => x"98ffc348",
    89 => x"66d07c70",
    90 => x"c329d049",
    91 => x"7c7199ff",
    92 => x"c84966d0",
    93 => x"99ffc329",
    94 => x"66d07c71",
    95 => x"99ffc349",
    96 => x"49727c71",
    97 => x"487129d0",
    98 => x"7098ffc3",
    99 => x"c94b6c7c",
   100 => x"c34dfff0",
   101 => x"d005abff",
   102 => x"7cffc387",
   103 => x"8dc14b6c",
   104 => x"c387c602",
   105 => x"f002abff",
   106 => x"fe487387",
   107 => x"c01e87c3",
   108 => x"48d4ff49",
   109 => x"c178ffc3",
   110 => x"b7c8c381",
   111 => x"87f104a9",
   112 => x"731e4f26",
   113 => x"c487e71e",
   114 => x"c04bdff8",
   115 => x"f0ffc01e",
   116 => x"fd49f7c1",
   117 => x"86c487e3",
   118 => x"c005a8c1",
   119 => x"d4ff87ea",
   120 => x"78ffc348",
   121 => x"c0c0c0c1",
   122 => x"c01ec0c0",
   123 => x"e9c1f0e1",
   124 => x"87c5fd49",
   125 => x"987086c4",
   126 => x"ff87ca05",
   127 => x"ffc348d4",
   128 => x"cb48c178",
   129 => x"87e6fe87",
   130 => x"fe058bc1",
   131 => x"48c087fd",
   132 => x"1e87e2fc",
   133 => x"d4ff1e73",
   134 => x"78ffc348",
   135 => x"1ec04bd3",
   136 => x"c1f0ffc0",
   137 => x"d0fc49c1",
   138 => x"7086c487",
   139 => x"87ca0598",
   140 => x"c348d4ff",
   141 => x"48c178ff",
   142 => x"f1fd87cb",
   143 => x"058bc187",
   144 => x"c087dbff",
   145 => x"87edfb48",
   146 => x"5c5b5e0e",
   147 => x"4cd4ff0e",
   148 => x"c687dbfd",
   149 => x"e1c01eea",
   150 => x"49c8c1f0",
   151 => x"c487dafb",
   152 => x"02a8c186",
   153 => x"eafe87c8",
   154 => x"c148c087",
   155 => x"d6fa87e2",
   156 => x"cf497087",
   157 => x"c699ffff",
   158 => x"c802a9ea",
   159 => x"87d3fe87",
   160 => x"cbc148c0",
   161 => x"7cffc387",
   162 => x"fc4bf1c0",
   163 => x"987087f4",
   164 => x"87ebc002",
   165 => x"ffc01ec0",
   166 => x"49fac1f0",
   167 => x"c487dafa",
   168 => x"05987086",
   169 => x"ffc387d9",
   170 => x"c3496c7c",
   171 => x"7c7c7cff",
   172 => x"99c0c17c",
   173 => x"c187c402",
   174 => x"c087d548",
   175 => x"c287d148",
   176 => x"87c405ab",
   177 => x"87c848c0",
   178 => x"fe058bc1",
   179 => x"48c087fd",
   180 => x"1e87e0f9",
   181 => x"dac21e73",
   182 => x"78c148e0",
   183 => x"d0ff4bc7",
   184 => x"fb78c248",
   185 => x"d0ff87c8",
   186 => x"c078c348",
   187 => x"d0e5c01e",
   188 => x"f949c0c1",
   189 => x"86c487c3",
   190 => x"c105a8c1",
   191 => x"abc24b87",
   192 => x"c087c505",
   193 => x"87f9c048",
   194 => x"ff058bc1",
   195 => x"f7fc87d0",
   196 => x"e4dac287",
   197 => x"05987058",
   198 => x"1ec187cd",
   199 => x"c1f0ffc0",
   200 => x"d4f849d0",
   201 => x"ff86c487",
   202 => x"ffc348d4",
   203 => x"87ddc478",
   204 => x"58e8dac2",
   205 => x"c248d0ff",
   206 => x"48d4ff78",
   207 => x"c178ffc3",
   208 => x"87f1f748",
   209 => x"5c5b5e0e",
   210 => x"4a710e5d",
   211 => x"ff4dffc3",
   212 => x"7c754cd4",
   213 => x"c448d0ff",
   214 => x"7c7578c3",
   215 => x"ffc01e72",
   216 => x"49d8c1f0",
   217 => x"c487d2f7",
   218 => x"02987086",
   219 => x"48c187c5",
   220 => x"7587eec0",
   221 => x"7cfec37c",
   222 => x"d41ec0c8",
   223 => x"f6f44966",
   224 => x"7586c487",
   225 => x"757c757c",
   226 => x"e0dad87c",
   227 => x"6c7c754b",
   228 => x"c187c505",
   229 => x"87f5058b",
   230 => x"d0ff7c75",
   231 => x"c078c248",
   232 => x"87cdf648",
   233 => x"5c5b5e0e",
   234 => x"4b710e5d",
   235 => x"eec54cc0",
   236 => x"ff4adfcd",
   237 => x"ffc348d4",
   238 => x"c3486878",
   239 => x"c005a8fe",
   240 => x"d4ff87fe",
   241 => x"029b734d",
   242 => x"66d087cc",
   243 => x"f449731e",
   244 => x"86c487cc",
   245 => x"d0ff87d6",
   246 => x"78d1c448",
   247 => x"d07dffc3",
   248 => x"88c14866",
   249 => x"7058a6d4",
   250 => x"87f00598",
   251 => x"c348d4ff",
   252 => x"737878ff",
   253 => x"87c5059b",
   254 => x"d048d0ff",
   255 => x"4c4ac178",
   256 => x"fe058ac1",
   257 => x"487487ed",
   258 => x"1e87e6f4",
   259 => x"4a711e73",
   260 => x"d4ff4bc0",
   261 => x"78ffc348",
   262 => x"c448d0ff",
   263 => x"d4ff78c3",
   264 => x"78ffc348",
   265 => x"ffc01e72",
   266 => x"49d1c1f0",
   267 => x"c487caf4",
   268 => x"05987086",
   269 => x"c0c887d2",
   270 => x"4966cc1e",
   271 => x"c487e5fd",
   272 => x"ff4b7086",
   273 => x"78c248d0",
   274 => x"e8f34873",
   275 => x"5b5e0e87",
   276 => x"c00e5d5c",
   277 => x"f0ffc01e",
   278 => x"f349c9c1",
   279 => x"1ed287db",
   280 => x"49e8dac2",
   281 => x"c887fdfc",
   282 => x"c14cc086",
   283 => x"acb7d284",
   284 => x"c287f804",
   285 => x"bf97e8da",
   286 => x"99c0c349",
   287 => x"05a9c0c1",
   288 => x"c287e7c0",
   289 => x"bf97efda",
   290 => x"c231d049",
   291 => x"bf97f0da",
   292 => x"7232c84a",
   293 => x"f1dac2b1",
   294 => x"b14abf97",
   295 => x"ffcf4c71",
   296 => x"c19cffff",
   297 => x"c134ca84",
   298 => x"dac287e7",
   299 => x"49bf97f1",
   300 => x"99c631c1",
   301 => x"97f2dac2",
   302 => x"b7c74abf",
   303 => x"c2b1722a",
   304 => x"bf97edda",
   305 => x"9dcf4d4a",
   306 => x"97eedac2",
   307 => x"9ac34abf",
   308 => x"dac232ca",
   309 => x"4bbf97ef",
   310 => x"b27333c2",
   311 => x"97f0dac2",
   312 => x"c0c34bbf",
   313 => x"2bb7c69b",
   314 => x"81c2b273",
   315 => x"307148c1",
   316 => x"48c14970",
   317 => x"4d703075",
   318 => x"84c14c72",
   319 => x"c0c89471",
   320 => x"cc06adb7",
   321 => x"b734c187",
   322 => x"b7c0c82d",
   323 => x"f4ff01ad",
   324 => x"f0487487",
   325 => x"5e0e87db",
   326 => x"0e5d5c5b",
   327 => x"e3c286f8",
   328 => x"78c048ce",
   329 => x"1ec6dbc2",
   330 => x"defb49c0",
   331 => x"7086c487",
   332 => x"87c50598",
   333 => x"c0c948c0",
   334 => x"c14dc087",
   335 => x"d9f2c07e",
   336 => x"dbc249bf",
   337 => x"c8714afc",
   338 => x"87ddec4b",
   339 => x"c2059870",
   340 => x"c07ec087",
   341 => x"49bfd5f2",
   342 => x"4ad8dcc2",
   343 => x"ec4bc871",
   344 => x"987087c7",
   345 => x"c087c205",
   346 => x"c0026e7e",
   347 => x"e2c287fd",
   348 => x"c24dbfcc",
   349 => x"bf9fc4e3",
   350 => x"d6c5487e",
   351 => x"c705a8ea",
   352 => x"cce2c287",
   353 => x"87ce4dbf",
   354 => x"e9ca486e",
   355 => x"c502a8d5",
   356 => x"c748c087",
   357 => x"dbc287e3",
   358 => x"49751ec6",
   359 => x"c487ecf9",
   360 => x"05987086",
   361 => x"48c087c5",
   362 => x"c087cec7",
   363 => x"49bfd5f2",
   364 => x"4ad8dcc2",
   365 => x"ea4bc871",
   366 => x"987087ef",
   367 => x"c287c805",
   368 => x"c148cee3",
   369 => x"c087da78",
   370 => x"49bfd9f2",
   371 => x"4afcdbc2",
   372 => x"ea4bc871",
   373 => x"987087d3",
   374 => x"87c5c002",
   375 => x"d8c648c0",
   376 => x"c4e3c287",
   377 => x"c149bf97",
   378 => x"c005a9d5",
   379 => x"e3c287cd",
   380 => x"49bf97c5",
   381 => x"02a9eac2",
   382 => x"c087c5c0",
   383 => x"87f9c548",
   384 => x"97c6dbc2",
   385 => x"c3487ebf",
   386 => x"c002a8e9",
   387 => x"486e87ce",
   388 => x"02a8ebc3",
   389 => x"c087c5c0",
   390 => x"87ddc548",
   391 => x"97d1dbc2",
   392 => x"059949bf",
   393 => x"c287ccc0",
   394 => x"bf97d2db",
   395 => x"02a9c249",
   396 => x"c087c5c0",
   397 => x"87c1c548",
   398 => x"97d3dbc2",
   399 => x"e3c248bf",
   400 => x"4c7058ca",
   401 => x"c288c148",
   402 => x"c258cee3",
   403 => x"bf97d4db",
   404 => x"c2817549",
   405 => x"bf97d5db",
   406 => x"7232c84a",
   407 => x"e7c27ea1",
   408 => x"786e48db",
   409 => x"97d6dbc2",
   410 => x"a6c848bf",
   411 => x"cee3c258",
   412 => x"cfc202bf",
   413 => x"d5f2c087",
   414 => x"dcc249bf",
   415 => x"c8714ad8",
   416 => x"87e5e74b",
   417 => x"c0029870",
   418 => x"48c087c5",
   419 => x"c287eac3",
   420 => x"4cbfc6e3",
   421 => x"5cefe7c2",
   422 => x"97ebdbc2",
   423 => x"31c849bf",
   424 => x"97eadbc2",
   425 => x"49a14abf",
   426 => x"97ecdbc2",
   427 => x"32d04abf",
   428 => x"c249a172",
   429 => x"bf97eddb",
   430 => x"7232d84a",
   431 => x"66c449a1",
   432 => x"dbe7c291",
   433 => x"e7c281bf",
   434 => x"dbc259e3",
   435 => x"4abf97f3",
   436 => x"dbc232c8",
   437 => x"4bbf97f2",
   438 => x"dbc24aa2",
   439 => x"4bbf97f4",
   440 => x"a27333d0",
   441 => x"f5dbc24a",
   442 => x"cf4bbf97",
   443 => x"7333d89b",
   444 => x"e7c24aa2",
   445 => x"8ac25ae7",
   446 => x"e7c29274",
   447 => x"a17248e7",
   448 => x"87c1c178",
   449 => x"97d8dbc2",
   450 => x"31c849bf",
   451 => x"97d7dbc2",
   452 => x"49a14abf",
   453 => x"ffc731c5",
   454 => x"c229c981",
   455 => x"c259efe7",
   456 => x"bf97dddb",
   457 => x"c232c84a",
   458 => x"bf97dcdb",
   459 => x"c44aa24b",
   460 => x"826e9266",
   461 => x"5aebe7c2",
   462 => x"48e3e7c2",
   463 => x"e7c278c0",
   464 => x"a17248df",
   465 => x"efe7c278",
   466 => x"e3e7c248",
   467 => x"e7c278bf",
   468 => x"e7c248f3",
   469 => x"c278bfe7",
   470 => x"02bfcee3",
   471 => x"7487c9c0",
   472 => x"7030c448",
   473 => x"87c9c07e",
   474 => x"bfebe7c2",
   475 => x"7030c448",
   476 => x"d2e3c27e",
   477 => x"c1786e48",
   478 => x"268ef848",
   479 => x"264c264d",
   480 => x"0e4f264b",
   481 => x"5d5c5b5e",
   482 => x"c24a710e",
   483 => x"02bfcee3",
   484 => x"4b7287cb",
   485 => x"4d722bc7",
   486 => x"c99dffc1",
   487 => x"c84b7287",
   488 => x"c34d722b",
   489 => x"e7c29dff",
   490 => x"c083bfdb",
   491 => x"abbfd1f2",
   492 => x"c087d902",
   493 => x"c25bd5f2",
   494 => x"731ec6db",
   495 => x"87cbf149",
   496 => x"987086c4",
   497 => x"c087c505",
   498 => x"87e6c048",
   499 => x"bfcee3c2",
   500 => x"7587d202",
   501 => x"c291c449",
   502 => x"6981c6db",
   503 => x"ffffcf4c",
   504 => x"cb9cffff",
   505 => x"c2497587",
   506 => x"c6dbc291",
   507 => x"4c699f81",
   508 => x"c6fe4874",
   509 => x"5b5e0e87",
   510 => x"f80e5d5c",
   511 => x"9c4c7186",
   512 => x"c087c505",
   513 => x"87c0c348",
   514 => x"487ea4c8",
   515 => x"66d878c0",
   516 => x"d887c702",
   517 => x"05bf9766",
   518 => x"48c087c5",
   519 => x"c087e9c2",
   520 => x"4949c11e",
   521 => x"c487d3ca",
   522 => x"9d4d7086",
   523 => x"87c2c102",
   524 => x"4ad6e3c2",
   525 => x"e04966d8",
   526 => x"987087d4",
   527 => x"87f2c002",
   528 => x"66d84a75",
   529 => x"e04bcb49",
   530 => x"987087f9",
   531 => x"87e2c002",
   532 => x"9d751ec0",
   533 => x"c887c702",
   534 => x"78c048a6",
   535 => x"a6c887c5",
   536 => x"c878c148",
   537 => x"d1c94966",
   538 => x"7086c487",
   539 => x"fe059d4d",
   540 => x"9d7587fe",
   541 => x"87cec102",
   542 => x"6e49a5dc",
   543 => x"da786948",
   544 => x"a6c449a5",
   545 => x"78a4c448",
   546 => x"c448699f",
   547 => x"c2780866",
   548 => x"02bfcee3",
   549 => x"a5d487d2",
   550 => x"49699f49",
   551 => x"99ffffc0",
   552 => x"30d04871",
   553 => x"87c27e70",
   554 => x"486e7ec0",
   555 => x"80bf66c4",
   556 => x"780866c4",
   557 => x"a4cc7cc0",
   558 => x"bf66c449",
   559 => x"49a4d079",
   560 => x"48c179c0",
   561 => x"48c087c2",
   562 => x"eefa8ef8",
   563 => x"5b5e0e87",
   564 => x"4c710e5c",
   565 => x"cbc1029c",
   566 => x"49a4c887",
   567 => x"c3c10269",
   568 => x"cc496c87",
   569 => x"80714866",
   570 => x"7058a6d0",
   571 => x"cae3c2b9",
   572 => x"baff4abf",
   573 => x"99719972",
   574 => x"87e5c002",
   575 => x"6b4ba4c4",
   576 => x"87fff949",
   577 => x"e3c27b70",
   578 => x"6c49bfc6",
   579 => x"cc7c7181",
   580 => x"e3c2b966",
   581 => x"ff4abfca",
   582 => x"719972ba",
   583 => x"dbff0599",
   584 => x"7c66cc87",
   585 => x"1e87d6f9",
   586 => x"4b711e73",
   587 => x"87c7029b",
   588 => x"6949a3c8",
   589 => x"c087c505",
   590 => x"87f6c048",
   591 => x"bfdfe7c2",
   592 => x"4aa3c449",
   593 => x"8ac24a6a",
   594 => x"bfc6e3c2",
   595 => x"49a17292",
   596 => x"bfcae3c2",
   597 => x"729a6b4a",
   598 => x"f2c049a1",
   599 => x"66c859d5",
   600 => x"e6ea711e",
   601 => x"7086c487",
   602 => x"87c40598",
   603 => x"87c248c0",
   604 => x"caf848c1",
   605 => x"1e731e87",
   606 => x"029b4b71",
   607 => x"a3c887c7",
   608 => x"c5056949",
   609 => x"c048c087",
   610 => x"e7c287f6",
   611 => x"c449bfdf",
   612 => x"4a6a4aa3",
   613 => x"e3c28ac2",
   614 => x"7292bfc6",
   615 => x"e3c249a1",
   616 => x"6b4abfca",
   617 => x"49a1729a",
   618 => x"59d5f2c0",
   619 => x"711e66c8",
   620 => x"c487d1e6",
   621 => x"05987086",
   622 => x"48c087c4",
   623 => x"48c187c2",
   624 => x"0e87fcf6",
   625 => x"5d5c5b5e",
   626 => x"4b711e0e",
   627 => x"734d66d4",
   628 => x"ccc1029b",
   629 => x"49a3c887",
   630 => x"c4c10269",
   631 => x"4ca3d087",
   632 => x"bfcae3c2",
   633 => x"6cb9ff49",
   634 => x"d47e994a",
   635 => x"cd06a966",
   636 => x"7c7bc087",
   637 => x"c44aa3cc",
   638 => x"796a49a3",
   639 => x"497287ca",
   640 => x"d499c0f8",
   641 => x"8d714d66",
   642 => x"29c94975",
   643 => x"49731e71",
   644 => x"c287fafa",
   645 => x"731ec6db",
   646 => x"87cbfc49",
   647 => x"66d486c8",
   648 => x"d6f5267c",
   649 => x"1e731e87",
   650 => x"029b4b71",
   651 => x"c287e4c0",
   652 => x"735bf3e7",
   653 => x"c28ac24a",
   654 => x"49bfc6e3",
   655 => x"dfe7c292",
   656 => x"807248bf",
   657 => x"58f7e7c2",
   658 => x"30c44871",
   659 => x"58d6e3c2",
   660 => x"c287edc0",
   661 => x"c248efe7",
   662 => x"78bfe3e7",
   663 => x"48f3e7c2",
   664 => x"bfe7e7c2",
   665 => x"cee3c278",
   666 => x"87c902bf",
   667 => x"bfc6e3c2",
   668 => x"c731c449",
   669 => x"ebe7c287",
   670 => x"31c449bf",
   671 => x"59d6e3c2",
   672 => x"0e87fcf3",
   673 => x"0e5c5b5e",
   674 => x"4bc04a71",
   675 => x"c0029a72",
   676 => x"a2da87e0",
   677 => x"4b699f49",
   678 => x"bfcee3c2",
   679 => x"d487cf02",
   680 => x"699f49a2",
   681 => x"ffc04c49",
   682 => x"34d09cff",
   683 => x"4cc087c2",
   684 => x"4973b374",
   685 => x"f387eefd",
   686 => x"5e0e87c3",
   687 => x"0e5d5c5b",
   688 => x"4a7186f4",
   689 => x"9a727ec0",
   690 => x"c287d802",
   691 => x"c048c2db",
   692 => x"fadac278",
   693 => x"f3e7c248",
   694 => x"dac278bf",
   695 => x"e7c248fe",
   696 => x"c278bfef",
   697 => x"c048e3e3",
   698 => x"d2e3c250",
   699 => x"dbc249bf",
   700 => x"714abfc2",
   701 => x"c9c403aa",
   702 => x"cf497287",
   703 => x"e9c00599",
   704 => x"d1f2c087",
   705 => x"fadac248",
   706 => x"dbc278bf",
   707 => x"dac21ec6",
   708 => x"c249bffa",
   709 => x"c148fada",
   710 => x"e37178a1",
   711 => x"86c487ed",
   712 => x"48cdf2c0",
   713 => x"78c6dbc2",
   714 => x"f2c087cc",
   715 => x"c048bfcd",
   716 => x"f2c080e0",
   717 => x"dbc258d1",
   718 => x"c148bfc2",
   719 => x"c6dbc280",
   720 => x"0c8d2758",
   721 => x"97bf0000",
   722 => x"029d4dbf",
   723 => x"c387e3c2",
   724 => x"c202ade5",
   725 => x"f2c087dc",
   726 => x"cb4bbfcd",
   727 => x"4c1149a3",
   728 => x"c105accf",
   729 => x"497587d2",
   730 => x"89c199df",
   731 => x"e3c291cd",
   732 => x"a3c181d6",
   733 => x"c351124a",
   734 => x"51124aa3",
   735 => x"124aa3c5",
   736 => x"4aa3c751",
   737 => x"a3c95112",
   738 => x"ce51124a",
   739 => x"51124aa3",
   740 => x"124aa3d0",
   741 => x"4aa3d251",
   742 => x"a3d45112",
   743 => x"d651124a",
   744 => x"51124aa3",
   745 => x"124aa3d8",
   746 => x"4aa3dc51",
   747 => x"a3de5112",
   748 => x"c151124a",
   749 => x"87fac07e",
   750 => x"99c84974",
   751 => x"87ebc005",
   752 => x"99d04974",
   753 => x"dc87d105",
   754 => x"cbc00266",
   755 => x"dc497387",
   756 => x"98700f66",
   757 => x"87d3c002",
   758 => x"c6c0056e",
   759 => x"d6e3c287",
   760 => x"c050c048",
   761 => x"48bfcdf2",
   762 => x"c287ddc2",
   763 => x"c048e3e3",
   764 => x"e3c27e50",
   765 => x"c249bfd2",
   766 => x"4abfc2db",
   767 => x"fb04aa71",
   768 => x"e7c287f7",
   769 => x"c005bff3",
   770 => x"e3c287c8",
   771 => x"c102bfce",
   772 => x"dac287f4",
   773 => x"ed49bffe",
   774 => x"dbc287e9",
   775 => x"a6c458c2",
   776 => x"fedac248",
   777 => x"e3c278bf",
   778 => x"c002bfce",
   779 => x"66c487d8",
   780 => x"ffffcf49",
   781 => x"a999f8ff",
   782 => x"87c5c002",
   783 => x"e1c04cc0",
   784 => x"c04cc187",
   785 => x"66c487dc",
   786 => x"f8ffcf49",
   787 => x"c002a999",
   788 => x"a6c887c8",
   789 => x"c078c048",
   790 => x"a6c887c5",
   791 => x"c878c148",
   792 => x"9c744c66",
   793 => x"87dec005",
   794 => x"c24966c4",
   795 => x"c6e3c289",
   796 => x"e7c291bf",
   797 => x"7148bfdf",
   798 => x"fedac280",
   799 => x"c2dbc258",
   800 => x"f978c048",
   801 => x"48c087e3",
   802 => x"eeeb8ef4",
   803 => x"00000087",
   804 => x"ffffff00",
   805 => x"000c9dff",
   806 => x"000ca600",
   807 => x"54414600",
   808 => x"20203233",
   809 => x"41460020",
   810 => x"20363154",
   811 => x"1e002020",
   812 => x"c348d4ff",
   813 => x"486878ff",
   814 => x"ff1e4f26",
   815 => x"ffc348d4",
   816 => x"48d0ff78",
   817 => x"ff78e1c0",
   818 => x"78d448d4",
   819 => x"48f7e7c2",
   820 => x"50bfd4ff",
   821 => x"ff1e4f26",
   822 => x"e0c048d0",
   823 => x"1e4f2678",
   824 => x"7087ccff",
   825 => x"c6029949",
   826 => x"a9fbc087",
   827 => x"7187f105",
   828 => x"0e4f2648",
   829 => x"0e5c5b5e",
   830 => x"4cc04b71",
   831 => x"7087f0fe",
   832 => x"c0029949",
   833 => x"ecc087f9",
   834 => x"f2c002a9",
   835 => x"a9fbc087",
   836 => x"87ebc002",
   837 => x"acb766cc",
   838 => x"d087c703",
   839 => x"87c20266",
   840 => x"99715371",
   841 => x"c187c202",
   842 => x"87c3fe84",
   843 => x"02994970",
   844 => x"ecc087cd",
   845 => x"87c702a9",
   846 => x"05a9fbc0",
   847 => x"d087d5ff",
   848 => x"87c30266",
   849 => x"c07b97c0",
   850 => x"c405a9ec",
   851 => x"c54a7487",
   852 => x"c04a7487",
   853 => x"48728a0a",
   854 => x"4d2687c2",
   855 => x"4b264c26",
   856 => x"fd1e4f26",
   857 => x"497087c9",
   858 => x"aaf0c04a",
   859 => x"c087c904",
   860 => x"c301aaf9",
   861 => x"8af0c087",
   862 => x"04aac1c1",
   863 => x"dac187c9",
   864 => x"87c301aa",
   865 => x"728af7c0",
   866 => x"0e4f2648",
   867 => x"5d5c5b5e",
   868 => x"7186f80e",
   869 => x"fc4dc04c",
   870 => x"4bc087e0",
   871 => x"97eaf8c0",
   872 => x"a9c049bf",
   873 => x"fc87cf04",
   874 => x"83c187f5",
   875 => x"97eaf8c0",
   876 => x"06ab49bf",
   877 => x"f8c087f1",
   878 => x"02bf97ea",
   879 => x"eefb87cf",
   880 => x"99497087",
   881 => x"c087c602",
   882 => x"f105a9ec",
   883 => x"fb4bc087",
   884 => x"7e7087dd",
   885 => x"c887d8fb",
   886 => x"d2fb58a6",
   887 => x"c14a7087",
   888 => x"49a4c883",
   889 => x"6e496997",
   890 => x"87da05a9",
   891 => x"9749a4c9",
   892 => x"66c44969",
   893 => x"87ce05a9",
   894 => x"9749a4ca",
   895 => x"05aa4969",
   896 => x"4dc187c4",
   897 => x"486e87d4",
   898 => x"02a8ecc0",
   899 => x"486e87c8",
   900 => x"05a8fbc0",
   901 => x"4bc087c4",
   902 => x"9d754dc1",
   903 => x"87effe02",
   904 => x"7387f3fa",
   905 => x"fc8ef848",
   906 => x"0e0087f0",
   907 => x"5d5c5b5e",
   908 => x"7186f80e",
   909 => x"4bd4ff7e",
   910 => x"e7c21e6e",
   911 => x"f4e649fc",
   912 => x"7086c487",
   913 => x"eac40298",
   914 => x"dae3c187",
   915 => x"496e4dbf",
   916 => x"c887f8fc",
   917 => x"987058a6",
   918 => x"c487c505",
   919 => x"78c148a6",
   920 => x"c548d0ff",
   921 => x"7bd5c178",
   922 => x"c14966c4",
   923 => x"c131c689",
   924 => x"bf97d8e3",
   925 => x"b071484a",
   926 => x"d0ff7b70",
   927 => x"c278c448",
   928 => x"bf97f7e7",
   929 => x"0299d049",
   930 => x"78c587d7",
   931 => x"c07bd6c1",
   932 => x"7bffc34a",
   933 => x"e0c082c1",
   934 => x"87f504aa",
   935 => x"c448d0ff",
   936 => x"7bffc378",
   937 => x"c548d0ff",
   938 => x"7bd3c178",
   939 => x"78c47bc1",
   940 => x"06adb7c0",
   941 => x"c287ebc2",
   942 => x"4cbfc4e8",
   943 => x"c2029c8d",
   944 => x"dbc287c2",
   945 => x"a6c47ec6",
   946 => x"78c0c848",
   947 => x"acb7c08c",
   948 => x"c887c603",
   949 => x"c078a4c0",
   950 => x"f7e7c24c",
   951 => x"d049bf97",
   952 => x"87d00299",
   953 => x"e7c21ec0",
   954 => x"fae849fc",
   955 => x"7086c487",
   956 => x"87f5c04a",
   957 => x"1ec6dbc2",
   958 => x"49fce7c2",
   959 => x"c487e8e8",
   960 => x"ff4a7086",
   961 => x"c5c848d0",
   962 => x"7bd4c178",
   963 => x"7bbf976e",
   964 => x"80c1486e",
   965 => x"66c47e70",
   966 => x"c888c148",
   967 => x"987058a6",
   968 => x"87e8ff05",
   969 => x"c448d0ff",
   970 => x"059a7278",
   971 => x"48c087c5",
   972 => x"c187c2c1",
   973 => x"fce7c21e",
   974 => x"87d1e649",
   975 => x"9c7486c4",
   976 => x"87fefd05",
   977 => x"06adb7c0",
   978 => x"e7c287d1",
   979 => x"78c048fc",
   980 => x"78c080d0",
   981 => x"e8c280f4",
   982 => x"c078bfc8",
   983 => x"fd01adb7",
   984 => x"d0ff87d5",
   985 => x"c178c548",
   986 => x"7bc07bd3",
   987 => x"48c178c4",
   988 => x"c087c2c0",
   989 => x"268ef848",
   990 => x"264c264d",
   991 => x"0e4f264b",
   992 => x"5d5c5b5e",
   993 => x"4b711e0e",
   994 => x"ab4d4cc0",
   995 => x"87e8c004",
   996 => x"1ecbf6c0",
   997 => x"c4029d75",
   998 => x"c24ac087",
   999 => x"724ac187",
  1000 => x"87d6ec49",
  1001 => x"7e7086c4",
  1002 => x"056e84c1",
  1003 => x"4c7387c2",
  1004 => x"ac7385c1",
  1005 => x"87d8ff06",
  1006 => x"fe26486e",
  1007 => x"5e0e87f9",
  1008 => x"710e5c5b",
  1009 => x"0266cc4b",
  1010 => x"c04c87d8",
  1011 => x"d8028cf0",
  1012 => x"c14a7487",
  1013 => x"87d1028a",
  1014 => x"87cd028a",
  1015 => x"87c9028a",
  1016 => x"497387d9",
  1017 => x"d287c4f9",
  1018 => x"c01e7487",
  1019 => x"f7d8c149",
  1020 => x"731e7487",
  1021 => x"efd8c149",
  1022 => x"fd86c887",
  1023 => x"5e0e87fb",
  1024 => x"0e5d5c5b",
  1025 => x"494c711e",
  1026 => x"e8c291de",
  1027 => x"85714de4",
  1028 => x"c1026d97",
  1029 => x"e8c287dc",
  1030 => x"7449bfd0",
  1031 => x"defd7181",
  1032 => x"487e7087",
  1033 => x"f2c00298",
  1034 => x"d8e8c287",
  1035 => x"cb4a704b",
  1036 => x"f2c1ff49",
  1037 => x"cb4b7487",
  1038 => x"ece3c193",
  1039 => x"c183c483",
  1040 => x"747bf6c1",
  1041 => x"d0c1c149",
  1042 => x"c17b7587",
  1043 => x"bf97d9e3",
  1044 => x"e8c21e49",
  1045 => x"e5fd49d8",
  1046 => x"7486c487",
  1047 => x"f8c0c149",
  1048 => x"c149c087",
  1049 => x"c287d7c2",
  1050 => x"c048f8e7",
  1051 => x"de49c178",
  1052 => x"fc2687cd",
  1053 => x"6f4c87c1",
  1054 => x"6e696461",
  1055 => x"2e2e2e67",
  1056 => x"1e731e00",
  1057 => x"c2494a71",
  1058 => x"81bfd0e8",
  1059 => x"87effb71",
  1060 => x"029b4b70",
  1061 => x"e74987c4",
  1062 => x"e8c287e9",
  1063 => x"78c048d0",
  1064 => x"dadd49c1",
  1065 => x"87d3fb87",
  1066 => x"c149c01e",
  1067 => x"2687cfc1",
  1068 => x"4a711e4f",
  1069 => x"c191cb49",
  1070 => x"c881ece3",
  1071 => x"c2481181",
  1072 => x"c258fce7",
  1073 => x"c048d0e8",
  1074 => x"dc49c178",
  1075 => x"4f2687f1",
  1076 => x"0299711e",
  1077 => x"e5c187d2",
  1078 => x"50c048c1",
  1079 => x"c2c180f7",
  1080 => x"e3c140f1",
  1081 => x"87ce78e5",
  1082 => x"48fde4c1",
  1083 => x"78dee3c1",
  1084 => x"c2c180fc",
  1085 => x"4f2678e8",
  1086 => x"5c5b5e0e",
  1087 => x"86f40e5d",
  1088 => x"4dc6dbc2",
  1089 => x"a6c44cc0",
  1090 => x"c278c048",
  1091 => x"48bfd0e8",
  1092 => x"c106a8c0",
  1093 => x"dbc287c0",
  1094 => x"029848c6",
  1095 => x"c087f7c0",
  1096 => x"c81ecbf6",
  1097 => x"87c70266",
  1098 => x"c048a6c4",
  1099 => x"c487c578",
  1100 => x"78c148a6",
  1101 => x"e64966c4",
  1102 => x"86c487c0",
  1103 => x"84c14d70",
  1104 => x"c14866c4",
  1105 => x"58a6c880",
  1106 => x"bfd0e8c2",
  1107 => x"87c603ac",
  1108 => x"ff059d75",
  1109 => x"4cc087c9",
  1110 => x"c3029d75",
  1111 => x"f6c087dc",
  1112 => x"66c81ecb",
  1113 => x"cc87c702",
  1114 => x"78c048a6",
  1115 => x"a6cc87c5",
  1116 => x"cc78c148",
  1117 => x"c1e54966",
  1118 => x"7086c487",
  1119 => x"0298487e",
  1120 => x"4987e4c2",
  1121 => x"699781cb",
  1122 => x"0299d049",
  1123 => x"7487d4c1",
  1124 => x"c191cb49",
  1125 => x"c181ece3",
  1126 => x"c879c1c2",
  1127 => x"51ffc381",
  1128 => x"91de4974",
  1129 => x"4de4e8c2",
  1130 => x"c1c28571",
  1131 => x"a5c17d97",
  1132 => x"51e0c049",
  1133 => x"97d6e3c2",
  1134 => x"87d202bf",
  1135 => x"a5c284c1",
  1136 => x"d6e3c24b",
  1137 => x"fe49db4a",
  1138 => x"c187dcfb",
  1139 => x"a5cd87d9",
  1140 => x"c151c049",
  1141 => x"4ba5c284",
  1142 => x"49cb4a6e",
  1143 => x"87c7fbfe",
  1144 => x"7487c4c1",
  1145 => x"c191cb49",
  1146 => x"c081ece3",
  1147 => x"c279feff",
  1148 => x"bf97d6e3",
  1149 => x"7487d802",
  1150 => x"c191de49",
  1151 => x"e4e8c284",
  1152 => x"c283714b",
  1153 => x"dd4ad6e3",
  1154 => x"dafafe49",
  1155 => x"7487d887",
  1156 => x"c293de4b",
  1157 => x"cb83e4e8",
  1158 => x"51c049a3",
  1159 => x"6e7384c1",
  1160 => x"fe49cb4a",
  1161 => x"c487c0fa",
  1162 => x"80c14866",
  1163 => x"c758a6c8",
  1164 => x"c5c003ac",
  1165 => x"fc056e87",
  1166 => x"487487e4",
  1167 => x"f6f48ef4",
  1168 => x"1e731e87",
  1169 => x"cb494b71",
  1170 => x"ece3c191",
  1171 => x"4aa1c881",
  1172 => x"48d8e3c1",
  1173 => x"a1c95012",
  1174 => x"eaf8c04a",
  1175 => x"ca501248",
  1176 => x"d9e3c181",
  1177 => x"c1501148",
  1178 => x"bf97d9e3",
  1179 => x"49c01e49",
  1180 => x"c287cbf5",
  1181 => x"de48f8e7",
  1182 => x"d649c178",
  1183 => x"f32687c1",
  1184 => x"5e0e87f9",
  1185 => x"0e5d5c5b",
  1186 => x"4d7186f4",
  1187 => x"c191cb49",
  1188 => x"c881ece3",
  1189 => x"a1ca4aa1",
  1190 => x"48a6c47e",
  1191 => x"bfc0ecc2",
  1192 => x"bf976e78",
  1193 => x"4866c44b",
  1194 => x"4b702873",
  1195 => x"cc48124c",
  1196 => x"9c7058a6",
  1197 => x"81c984c1",
  1198 => x"b7496997",
  1199 => x"87c204ac",
  1200 => x"976e4cc0",
  1201 => x"66c84abf",
  1202 => x"ff317249",
  1203 => x"9966c4b9",
  1204 => x"30724874",
  1205 => x"71484a70",
  1206 => x"c4ecc2b0",
  1207 => x"f8e4c058",
  1208 => x"d449c087",
  1209 => x"497587d9",
  1210 => x"87edf6c0",
  1211 => x"c6f28ef4",
  1212 => x"1e731e87",
  1213 => x"fe494b71",
  1214 => x"497387c8",
  1215 => x"f187c3fe",
  1216 => x"731e87f9",
  1217 => x"c64b711e",
  1218 => x"c0024aa3",
  1219 => x"8ac187e3",
  1220 => x"8a87d602",
  1221 => x"87e8c102",
  1222 => x"cac1028a",
  1223 => x"c0028a87",
  1224 => x"028a87ef",
  1225 => x"e9c187d9",
  1226 => x"f649c787",
  1227 => x"ecc187c3",
  1228 => x"f8e7c287",
  1229 => x"c178df48",
  1230 => x"87c3d349",
  1231 => x"c287dec1",
  1232 => x"02bfd0e8",
  1233 => x"4887cbc1",
  1234 => x"e8c288c1",
  1235 => x"c1c158d4",
  1236 => x"d4e8c287",
  1237 => x"f9c002bf",
  1238 => x"d0e8c287",
  1239 => x"80c148bf",
  1240 => x"58d4e8c2",
  1241 => x"c287ebc0",
  1242 => x"49bfd0e8",
  1243 => x"e8c289c6",
  1244 => x"b7c059d4",
  1245 => x"87da03a9",
  1246 => x"48d0e8c2",
  1247 => x"87d278c0",
  1248 => x"bfd4e8c2",
  1249 => x"c287cb02",
  1250 => x"48bfd0e8",
  1251 => x"e8c280c6",
  1252 => x"49c058d4",
  1253 => x"7387e8d1",
  1254 => x"fcf3c049",
  1255 => x"87dbef87",
  1256 => x"5c5b5e0e",
  1257 => x"d4ff0e5d",
  1258 => x"59a6dc86",
  1259 => x"c048a6c8",
  1260 => x"c180c478",
  1261 => x"c47866c0",
  1262 => x"c478c180",
  1263 => x"c278c180",
  1264 => x"c148d4e8",
  1265 => x"f8e7c278",
  1266 => x"a8de48bf",
  1267 => x"f487c905",
  1268 => x"a6cc87e6",
  1269 => x"87e6cf58",
  1270 => x"e487dfe3",
  1271 => x"cee387c1",
  1272 => x"c04c7087",
  1273 => x"c102acfb",
  1274 => x"66d887fb",
  1275 => x"87edc105",
  1276 => x"4a66fcc0",
  1277 => x"7e6a82c4",
  1278 => x"dfc11e72",
  1279 => x"66c448f3",
  1280 => x"4aa1c849",
  1281 => x"aa714120",
  1282 => x"1087f905",
  1283 => x"c04a2651",
  1284 => x"c14866fc",
  1285 => x"6a78c1c9",
  1286 => x"7481c749",
  1287 => x"66fcc051",
  1288 => x"c181c849",
  1289 => x"66fcc051",
  1290 => x"c081c949",
  1291 => x"66fcc051",
  1292 => x"c081ca49",
  1293 => x"d81ec151",
  1294 => x"c8496a1e",
  1295 => x"87f3e281",
  1296 => x"c0c186c8",
  1297 => x"a8c04866",
  1298 => x"c887c701",
  1299 => x"78c148a6",
  1300 => x"c0c187ce",
  1301 => x"88c14866",
  1302 => x"c358a6d0",
  1303 => x"87ffe187",
  1304 => x"c248a6d0",
  1305 => x"029c7478",
  1306 => x"c887cfcd",
  1307 => x"c4c14866",
  1308 => x"cd03a866",
  1309 => x"a6dc87c4",
  1310 => x"e878c048",
  1311 => x"e078c080",
  1312 => x"4c7087ed",
  1313 => x"05acd0c1",
  1314 => x"c487d7c2",
  1315 => x"d1e37e66",
  1316 => x"58a6c887",
  1317 => x"7087d8e0",
  1318 => x"acecc04c",
  1319 => x"87edc105",
  1320 => x"cb4966c8",
  1321 => x"66fcc091",
  1322 => x"4aa1c481",
  1323 => x"a1c84d6a",
  1324 => x"5266c44a",
  1325 => x"79f1c2c1",
  1326 => x"87f3dfff",
  1327 => x"029c4c70",
  1328 => x"fbc087d9",
  1329 => x"87d302ac",
  1330 => x"dfff5574",
  1331 => x"4c7087e1",
  1332 => x"87c7029c",
  1333 => x"05acfbc0",
  1334 => x"c087edff",
  1335 => x"c1c255e0",
  1336 => x"7d97c055",
  1337 => x"6e4866d8",
  1338 => x"87db05a8",
  1339 => x"cc4866c8",
  1340 => x"ca04a866",
  1341 => x"4866c887",
  1342 => x"a6cc80c1",
  1343 => x"cc87c858",
  1344 => x"88c14866",
  1345 => x"ff58a6d0",
  1346 => x"7087e4de",
  1347 => x"acd0c14c",
  1348 => x"d487c805",
  1349 => x"80c14866",
  1350 => x"c158a6d8",
  1351 => x"fd02acd0",
  1352 => x"66c487e9",
  1353 => x"a866d848",
  1354 => x"87e0c905",
  1355 => x"48a6e0c0",
  1356 => x"487478c0",
  1357 => x"7088fbc0",
  1358 => x"0298487e",
  1359 => x"4887e2c9",
  1360 => x"7e7088cb",
  1361 => x"c1029848",
  1362 => x"c94887cd",
  1363 => x"487e7088",
  1364 => x"fec30298",
  1365 => x"88c44887",
  1366 => x"98487e70",
  1367 => x"4887ce02",
  1368 => x"7e7088c1",
  1369 => x"c3029848",
  1370 => x"d6c887e9",
  1371 => x"48a6dc87",
  1372 => x"ff78f0c0",
  1373 => x"7087f8dc",
  1374 => x"acecc04c",
  1375 => x"87c4c002",
  1376 => x"5ca6e0c0",
  1377 => x"02acecc0",
  1378 => x"dcff87cd",
  1379 => x"4c7087e1",
  1380 => x"05acecc0",
  1381 => x"c087f3ff",
  1382 => x"c002acec",
  1383 => x"dcff87c4",
  1384 => x"1ec087cd",
  1385 => x"66d01eca",
  1386 => x"c191cb49",
  1387 => x"714866c4",
  1388 => x"58a6cc80",
  1389 => x"c44866c8",
  1390 => x"58a6d080",
  1391 => x"49bf66cc",
  1392 => x"87efdcff",
  1393 => x"1ede1ec1",
  1394 => x"49bf66d4",
  1395 => x"87e3dcff",
  1396 => x"497086d0",
  1397 => x"8808c048",
  1398 => x"58a6e8c0",
  1399 => x"c006a8c0",
  1400 => x"e4c087ee",
  1401 => x"a8dd4866",
  1402 => x"87e4c003",
  1403 => x"49bf66c4",
  1404 => x"8166e4c0",
  1405 => x"c051e0c0",
  1406 => x"c14966e4",
  1407 => x"bf66c481",
  1408 => x"51c1c281",
  1409 => x"4966e4c0",
  1410 => x"66c481c2",
  1411 => x"51c081bf",
  1412 => x"c9c1486e",
  1413 => x"496e78c1",
  1414 => x"66d081c8",
  1415 => x"c9496e51",
  1416 => x"5166d481",
  1417 => x"81ca496e",
  1418 => x"d05166dc",
  1419 => x"80c14866",
  1420 => x"c858a6d4",
  1421 => x"66cc4866",
  1422 => x"cbc004a8",
  1423 => x"4866c887",
  1424 => x"a6cc80c1",
  1425 => x"87d9c558",
  1426 => x"c14866cc",
  1427 => x"58a6d088",
  1428 => x"ff87cec5",
  1429 => x"c087cbdc",
  1430 => x"ff58a6e8",
  1431 => x"c087c3dc",
  1432 => x"c058a6e0",
  1433 => x"c005a8ec",
  1434 => x"a6dc87ca",
  1435 => x"66e4c048",
  1436 => x"87c4c078",
  1437 => x"87f7d8ff",
  1438 => x"cb4966c8",
  1439 => x"66fcc091",
  1440 => x"70807148",
  1441 => x"82c84a7e",
  1442 => x"81ca496e",
  1443 => x"5166e4c0",
  1444 => x"c14966dc",
  1445 => x"66e4c081",
  1446 => x"7148c189",
  1447 => x"c1497030",
  1448 => x"7a977189",
  1449 => x"bfc0ecc2",
  1450 => x"66e4c049",
  1451 => x"4a6a9729",
  1452 => x"c0987148",
  1453 => x"6e58a6ec",
  1454 => x"6981c449",
  1455 => x"4866d84d",
  1456 => x"02a866c4",
  1457 => x"c487c8c0",
  1458 => x"78c048a6",
  1459 => x"c487c5c0",
  1460 => x"78c148a6",
  1461 => x"c01e66c4",
  1462 => x"49751ee0",
  1463 => x"87d3d8ff",
  1464 => x"4c7086c8",
  1465 => x"06acb7c0",
  1466 => x"7487d4c1",
  1467 => x"49e0c085",
  1468 => x"4b758974",
  1469 => x"4afcdfc1",
  1470 => x"eae6fe71",
  1471 => x"c085c287",
  1472 => x"c14866e0",
  1473 => x"a6e4c080",
  1474 => x"66e8c058",
  1475 => x"7081c149",
  1476 => x"c8c002a9",
  1477 => x"48a6c487",
  1478 => x"c5c078c0",
  1479 => x"48a6c487",
  1480 => x"66c478c1",
  1481 => x"49a4c21e",
  1482 => x"7148e0c0",
  1483 => x"1e497088",
  1484 => x"d6ff4975",
  1485 => x"86c887fd",
  1486 => x"01a8b7c0",
  1487 => x"c087c0ff",
  1488 => x"c00266e0",
  1489 => x"496e87d1",
  1490 => x"e0c081c9",
  1491 => x"486e5166",
  1492 => x"78c2cac1",
  1493 => x"6e87ccc0",
  1494 => x"c281c949",
  1495 => x"c1486e51",
  1496 => x"c878f1cb",
  1497 => x"66cc4866",
  1498 => x"cbc004a8",
  1499 => x"4866c887",
  1500 => x"a6cc80c1",
  1501 => x"87e9c058",
  1502 => x"c14866cc",
  1503 => x"58a6d088",
  1504 => x"ff87dec0",
  1505 => x"7087d8d5",
  1506 => x"87d5c04c",
  1507 => x"05acc6c1",
  1508 => x"d087c8c0",
  1509 => x"80c14866",
  1510 => x"ff58a6d4",
  1511 => x"7087c0d5",
  1512 => x"4866d44c",
  1513 => x"a6d880c1",
  1514 => x"029c7458",
  1515 => x"c887cbc0",
  1516 => x"c4c14866",
  1517 => x"f204a866",
  1518 => x"d4ff87fc",
  1519 => x"66c887d8",
  1520 => x"03a8c748",
  1521 => x"c287e5c0",
  1522 => x"c048d4e8",
  1523 => x"4966c878",
  1524 => x"fcc091cb",
  1525 => x"a1c48166",
  1526 => x"c04a6a4a",
  1527 => x"66c87952",
  1528 => x"cc80c148",
  1529 => x"a8c758a6",
  1530 => x"87dbff04",
  1531 => x"ff8ed4ff",
  1532 => x"4c87c4de",
  1533 => x"2064616f",
  1534 => x"00202e2a",
  1535 => x"1e00203a",
  1536 => x"4b711e73",
  1537 => x"87c6029b",
  1538 => x"48d0e8c2",
  1539 => x"1ec778c0",
  1540 => x"bfd0e8c2",
  1541 => x"ece3c11e",
  1542 => x"f8e7c21e",
  1543 => x"ffed49bf",
  1544 => x"c286cc87",
  1545 => x"49bff8e7",
  1546 => x"7387e5e2",
  1547 => x"87c8029b",
  1548 => x"49ece3c1",
  1549 => x"87f3e2c0",
  1550 => x"87ffdcff",
  1551 => x"d8e3c11e",
  1552 => x"c150c048",
  1553 => x"49bfcfe5",
  1554 => x"87dfd7ff",
  1555 => x"4f2648c0",
  1556 => x"87dfc71e",
  1557 => x"e6fe49c1",
  1558 => x"f6e9fe87",
  1559 => x"02987087",
  1560 => x"f2fe87cd",
  1561 => x"987087f0",
  1562 => x"c187c402",
  1563 => x"c087c24a",
  1564 => x"059a724a",
  1565 => x"1ec087ce",
  1566 => x"49ebe2c1",
  1567 => x"87deefc0",
  1568 => x"87fe86c4",
  1569 => x"48d0e8c2",
  1570 => x"e7c278c0",
  1571 => x"78c048f8",
  1572 => x"f6e2c11e",
  1573 => x"c5efc049",
  1574 => x"fe1ec087",
  1575 => x"497087de",
  1576 => x"87faeec0",
  1577 => x"f887cbc3",
  1578 => x"534f268e",
  1579 => x"61662044",
  1580 => x"64656c69",
  1581 => x"6f42002e",
  1582 => x"6e69746f",
  1583 => x"2e2e2e67",
  1584 => x"e2c01e00",
  1585 => x"f2c087e2",
  1586 => x"87f687ce",
  1587 => x"fd1e4f26",
  1588 => x"87ed87fe",
  1589 => x"4f2648c0",
  1590 => x"00010000",
  1591 => x"20800000",
  1592 => x"74697845",
  1593 => x"42208000",
  1594 => x"006b6361",
  1595 => x"00000ffe",
  1596 => x"00002a24",
  1597 => x"fe000000",
  1598 => x"4200000f",
  1599 => x"0000002a",
  1600 => x"0ffe0000",
  1601 => x"2a600000",
  1602 => x"00000000",
  1603 => x"000ffe00",
  1604 => x"002a7e00",
  1605 => x"00000000",
  1606 => x"00000ffe",
  1607 => x"00002a9c",
  1608 => x"fe000000",
  1609 => x"ba00000f",
  1610 => x"0000002a",
  1611 => x"0ffe0000",
  1612 => x"2ad80000",
  1613 => x"00000000",
  1614 => x"0010b100",
  1615 => x"00000000",
  1616 => x"00000000",
  1617 => x"00001302",
  1618 => x"00000000",
  1619 => x"53000000",
  1620 => x"42000019",
  1621 => x"20544f4f",
  1622 => x"52202020",
  1623 => x"1e004d4f",
  1624 => x"c048f0fe",
  1625 => x"7909cd78",
  1626 => x"1e4f2609",
  1627 => x"48bff0fe",
  1628 => x"fe1e4f26",
  1629 => x"78c148f0",
  1630 => x"fe1e4f26",
  1631 => x"78c048f0",
  1632 => x"711e4f26",
  1633 => x"5152c04a",
  1634 => x"5e0e4f26",
  1635 => x"0e5d5c5b",
  1636 => x"4d7186f4",
  1637 => x"c17e6d97",
  1638 => x"6c974ca5",
  1639 => x"58a6c848",
  1640 => x"66c4486e",
  1641 => x"87c505a8",
  1642 => x"e6c048ff",
  1643 => x"87caff87",
  1644 => x"9749a5c2",
  1645 => x"a3714b6c",
  1646 => x"4b6b974b",
  1647 => x"6e7e6c97",
  1648 => x"c880c148",
  1649 => x"98c758a6",
  1650 => x"7058a6cc",
  1651 => x"e1fe7c97",
  1652 => x"f4487387",
  1653 => x"264d268e",
  1654 => x"264b264c",
  1655 => x"5b5e0e4f",
  1656 => x"86f40e5c",
  1657 => x"66d84c71",
  1658 => x"9affc34a",
  1659 => x"974ba4c2",
  1660 => x"a173496c",
  1661 => x"97517249",
  1662 => x"486e7e6c",
  1663 => x"a6c880c1",
  1664 => x"cc98c758",
  1665 => x"547058a6",
  1666 => x"caff8ef4",
  1667 => x"fd1e1e87",
  1668 => x"bfe087e8",
  1669 => x"e0c0494a",
  1670 => x"cb0299c0",
  1671 => x"c21e7287",
  1672 => x"fe49f6eb",
  1673 => x"86c487f7",
  1674 => x"7087c0fd",
  1675 => x"87c2fd7e",
  1676 => x"1e4f2626",
  1677 => x"49f6ebc2",
  1678 => x"c187c7fd",
  1679 => x"fc49cde8",
  1680 => x"eec387dd",
  1681 => x"0e4f2687",
  1682 => x"5d5c5b5e",
  1683 => x"c24d710e",
  1684 => x"fc49f6eb",
  1685 => x"4b7087f4",
  1686 => x"04abb7c0",
  1687 => x"c387c2c3",
  1688 => x"c905abf0",
  1689 => x"ebecc187",
  1690 => x"c278c148",
  1691 => x"e0c387e3",
  1692 => x"87c905ab",
  1693 => x"48efecc1",
  1694 => x"d4c278c1",
  1695 => x"efecc187",
  1696 => x"87c602bf",
  1697 => x"4ca3c0c2",
  1698 => x"4c7387c2",
  1699 => x"bfebecc1",
  1700 => x"87e0c002",
  1701 => x"b7c44974",
  1702 => x"eec19129",
  1703 => x"4a7481c2",
  1704 => x"92c29acf",
  1705 => x"307248c1",
  1706 => x"baff4a70",
  1707 => x"98694872",
  1708 => x"87db7970",
  1709 => x"b7c44974",
  1710 => x"eec19129",
  1711 => x"4a7481c2",
  1712 => x"92c29acf",
  1713 => x"307248c3",
  1714 => x"69484a70",
  1715 => x"757970b0",
  1716 => x"f0c0059d",
  1717 => x"48d0ff87",
  1718 => x"ff78e1c8",
  1719 => x"78c548d4",
  1720 => x"bfefecc1",
  1721 => x"c387c302",
  1722 => x"ecc178e0",
  1723 => x"c602bfeb",
  1724 => x"48d4ff87",
  1725 => x"ff78f0c3",
  1726 => x"0b7b0bd4",
  1727 => x"c848d0ff",
  1728 => x"e0c078e1",
  1729 => x"efecc178",
  1730 => x"c178c048",
  1731 => x"c048ebec",
  1732 => x"f6ebc278",
  1733 => x"87f2f949",
  1734 => x"b7c04b70",
  1735 => x"fefc03ab",
  1736 => x"2648c087",
  1737 => x"264c264d",
  1738 => x"004f264b",
  1739 => x"00000000",
  1740 => x"1e000000",
  1741 => x"49724ac0",
  1742 => x"eec191c4",
  1743 => x"79c081c2",
  1744 => x"b7d082c1",
  1745 => x"87ee04aa",
  1746 => x"5e0e4f26",
  1747 => x"0e5d5c5b",
  1748 => x"e5f84d71",
  1749 => x"c44a7587",
  1750 => x"c1922ab7",
  1751 => x"7582c2ee",
  1752 => x"c29ccf4c",
  1753 => x"4b496a94",
  1754 => x"9bc32b74",
  1755 => x"307448c2",
  1756 => x"bcff4c70",
  1757 => x"98714874",
  1758 => x"f5f77a70",
  1759 => x"fe487387",
  1760 => x"000087e1",
  1761 => x"00000000",
  1762 => x"00000000",
  1763 => x"00000000",
  1764 => x"00000000",
  1765 => x"00000000",
  1766 => x"00000000",
  1767 => x"00000000",
  1768 => x"00000000",
  1769 => x"00000000",
  1770 => x"00000000",
  1771 => x"00000000",
  1772 => x"00000000",
  1773 => x"00000000",
  1774 => x"00000000",
  1775 => x"00000000",
  1776 => x"ff1e0000",
  1777 => x"e1c848d0",
  1778 => x"ff487178",
  1779 => x"267808d4",
  1780 => x"d0ff1e4f",
  1781 => x"78e1c848",
  1782 => x"d4ff4871",
  1783 => x"66c47808",
  1784 => x"08d4ff48",
  1785 => x"1e4f2678",
  1786 => x"66c44a71",
  1787 => x"49721e49",
  1788 => x"ff87deff",
  1789 => x"e0c048d0",
  1790 => x"4f262678",
  1791 => x"711e731e",
  1792 => x"4966c84b",
  1793 => x"c14a731e",
  1794 => x"ff49a2e0",
  1795 => x"c42687d9",
  1796 => x"264d2687",
  1797 => x"264b264c",
  1798 => x"d4ff1e4f",
  1799 => x"7affc34a",
  1800 => x"c048d0ff",
  1801 => x"7ade78e1",
  1802 => x"bfc0ecc2",
  1803 => x"c848497a",
  1804 => x"717a7028",
  1805 => x"7028d048",
  1806 => x"d848717a",
  1807 => x"ff7a7028",
  1808 => x"e0c048d0",
  1809 => x"1e4f2678",
  1810 => x"c848d0ff",
  1811 => x"487178c9",
  1812 => x"7808d4ff",
  1813 => x"711e4f26",
  1814 => x"87eb494a",
  1815 => x"c848d0ff",
  1816 => x"1e4f2678",
  1817 => x"4b711e73",
  1818 => x"bfd0ecc2",
  1819 => x"c287c302",
  1820 => x"d0ff87eb",
  1821 => x"78c9c848",
  1822 => x"e0c04873",
  1823 => x"08d4ffb0",
  1824 => x"c4ecc278",
  1825 => x"c878c048",
  1826 => x"87c50266",
  1827 => x"c249ffc3",
  1828 => x"c249c087",
  1829 => x"cc59ccec",
  1830 => x"87c60266",
  1831 => x"4ad5d5c5",
  1832 => x"ffcf87c4",
  1833 => x"ecc24aff",
  1834 => x"ecc25ad0",
  1835 => x"78c148d0",
  1836 => x"4d2687c4",
  1837 => x"4b264c26",
  1838 => x"5e0e4f26",
  1839 => x"0e5d5c5b",
  1840 => x"ecc24a71",
  1841 => x"724cbfcc",
  1842 => x"87cb029a",
  1843 => x"c191c849",
  1844 => x"714bd9f1",
  1845 => x"c187c483",
  1846 => x"c04bd9f5",
  1847 => x"7449134d",
  1848 => x"c8ecc299",
  1849 => x"b87148bf",
  1850 => x"7808d4ff",
  1851 => x"852cb7c1",
  1852 => x"04adb7c8",
  1853 => x"ecc287e7",
  1854 => x"c848bfc4",
  1855 => x"c8ecc280",
  1856 => x"87eefe58",
  1857 => x"711e731e",
  1858 => x"9a4a134b",
  1859 => x"7287cb02",
  1860 => x"87e6fe49",
  1861 => x"059a4a13",
  1862 => x"d9fe87f5",
  1863 => x"ecc21e87",
  1864 => x"c249bfc4",
  1865 => x"c148c4ec",
  1866 => x"c0c478a1",
  1867 => x"db03a9b7",
  1868 => x"48d4ff87",
  1869 => x"bfc8ecc2",
  1870 => x"c4ecc278",
  1871 => x"ecc249bf",
  1872 => x"a1c148c4",
  1873 => x"b7c0c478",
  1874 => x"87e504a9",
  1875 => x"c848d0ff",
  1876 => x"d0ecc278",
  1877 => x"2678c048",
  1878 => x"0000004f",
  1879 => x"00000000",
  1880 => x"00000000",
  1881 => x"00005f5f",
  1882 => x"03030000",
  1883 => x"00030300",
  1884 => x"7f7f1400",
  1885 => x"147f7f14",
  1886 => x"2e240000",
  1887 => x"123a6b6b",
  1888 => x"366a4c00",
  1889 => x"32566c18",
  1890 => x"4f7e3000",
  1891 => x"683a7759",
  1892 => x"04000040",
  1893 => x"00000307",
  1894 => x"1c000000",
  1895 => x"0041633e",
  1896 => x"41000000",
  1897 => x"001c3e63",
  1898 => x"3e2a0800",
  1899 => x"2a3e1c1c",
  1900 => x"08080008",
  1901 => x"08083e3e",
  1902 => x"80000000",
  1903 => x"000060e0",
  1904 => x"08080000",
  1905 => x"08080808",
  1906 => x"00000000",
  1907 => x"00006060",
  1908 => x"30604000",
  1909 => x"03060c18",
  1910 => x"7f3e0001",
  1911 => x"3e7f4d59",
  1912 => x"06040000",
  1913 => x"00007f7f",
  1914 => x"63420000",
  1915 => x"464f5971",
  1916 => x"63220000",
  1917 => x"367f4949",
  1918 => x"161c1800",
  1919 => x"107f7f13",
  1920 => x"67270000",
  1921 => x"397d4545",
  1922 => x"7e3c0000",
  1923 => x"3079494b",
  1924 => x"01010000",
  1925 => x"070f7971",
  1926 => x"7f360000",
  1927 => x"367f4949",
  1928 => x"4f060000",
  1929 => x"1e3f6949",
  1930 => x"00000000",
  1931 => x"00006666",
  1932 => x"80000000",
  1933 => x"000066e6",
  1934 => x"08080000",
  1935 => x"22221414",
  1936 => x"14140000",
  1937 => x"14141414",
  1938 => x"22220000",
  1939 => x"08081414",
  1940 => x"03020000",
  1941 => x"060f5951",
  1942 => x"417f3e00",
  1943 => x"1e1f555d",
  1944 => x"7f7e0000",
  1945 => x"7e7f0909",
  1946 => x"7f7f0000",
  1947 => x"367f4949",
  1948 => x"3e1c0000",
  1949 => x"41414163",
  1950 => x"7f7f0000",
  1951 => x"1c3e6341",
  1952 => x"7f7f0000",
  1953 => x"41414949",
  1954 => x"7f7f0000",
  1955 => x"01010909",
  1956 => x"7f3e0000",
  1957 => x"7a7b4941",
  1958 => x"7f7f0000",
  1959 => x"7f7f0808",
  1960 => x"41000000",
  1961 => x"00417f7f",
  1962 => x"60200000",
  1963 => x"3f7f4040",
  1964 => x"087f7f00",
  1965 => x"4163361c",
  1966 => x"7f7f0000",
  1967 => x"40404040",
  1968 => x"067f7f00",
  1969 => x"7f7f060c",
  1970 => x"067f7f00",
  1971 => x"7f7f180c",
  1972 => x"7f3e0000",
  1973 => x"3e7f4141",
  1974 => x"7f7f0000",
  1975 => x"060f0909",
  1976 => x"417f3e00",
  1977 => x"407e7f61",
  1978 => x"7f7f0000",
  1979 => x"667f1909",
  1980 => x"6f260000",
  1981 => x"327b594d",
  1982 => x"01010000",
  1983 => x"01017f7f",
  1984 => x"7f3f0000",
  1985 => x"3f7f4040",
  1986 => x"3f0f0000",
  1987 => x"0f3f7070",
  1988 => x"307f7f00",
  1989 => x"7f7f3018",
  1990 => x"36634100",
  1991 => x"63361c1c",
  1992 => x"06030141",
  1993 => x"03067c7c",
  1994 => x"59716101",
  1995 => x"4143474d",
  1996 => x"7f000000",
  1997 => x"0041417f",
  1998 => x"06030100",
  1999 => x"6030180c",
  2000 => x"41000040",
  2001 => x"007f7f41",
  2002 => x"060c0800",
  2003 => x"080c0603",
  2004 => x"80808000",
  2005 => x"80808080",
  2006 => x"00000000",
  2007 => x"00040703",
  2008 => x"74200000",
  2009 => x"787c5454",
  2010 => x"7f7f0000",
  2011 => x"387c4444",
  2012 => x"7c380000",
  2013 => x"00444444",
  2014 => x"7c380000",
  2015 => x"7f7f4444",
  2016 => x"7c380000",
  2017 => x"185c5454",
  2018 => x"7e040000",
  2019 => x"0005057f",
  2020 => x"bc180000",
  2021 => x"7cfca4a4",
  2022 => x"7f7f0000",
  2023 => x"787c0404",
  2024 => x"00000000",
  2025 => x"00407d3d",
  2026 => x"80800000",
  2027 => x"007dfd80",
  2028 => x"7f7f0000",
  2029 => x"446c3810",
  2030 => x"00000000",
  2031 => x"00407f3f",
  2032 => x"0c7c7c00",
  2033 => x"787c0c18",
  2034 => x"7c7c0000",
  2035 => x"787c0404",
  2036 => x"7c380000",
  2037 => x"387c4444",
  2038 => x"fcfc0000",
  2039 => x"183c2424",
  2040 => x"3c180000",
  2041 => x"fcfc2424",
  2042 => x"7c7c0000",
  2043 => x"080c0404",
  2044 => x"5c480000",
  2045 => x"20745454",
  2046 => x"3f040000",
  2047 => x"0044447f",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
