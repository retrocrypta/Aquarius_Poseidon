
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom2 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"7c",x"3c",x"00",x"00"),
     1 => (x"7c",x"7c",x"40",x"40"),
     2 => (x"3c",x"1c",x"00",x"00"),
     3 => (x"1c",x"3c",x"60",x"60"),
     4 => (x"60",x"7c",x"3c",x"00"),
     5 => (x"3c",x"7c",x"60",x"30"),
     6 => (x"38",x"6c",x"44",x"00"),
     7 => (x"44",x"6c",x"38",x"10"),
     8 => (x"bc",x"1c",x"00",x"00"),
     9 => (x"1c",x"3c",x"60",x"e0"),
    10 => (x"64",x"44",x"00",x"00"),
    11 => (x"44",x"4c",x"5c",x"74"),
    12 => (x"08",x"08",x"00",x"00"),
    13 => (x"41",x"41",x"77",x"3e"),
    14 => (x"00",x"00",x"00",x"00"),
    15 => (x"00",x"00",x"7f",x"7f"),
    16 => (x"41",x"41",x"00",x"00"),
    17 => (x"08",x"08",x"3e",x"77"),
    18 => (x"01",x"01",x"02",x"00"),
    19 => (x"01",x"02",x"02",x"03"),
    20 => (x"7f",x"7f",x"7f",x"00"),
    21 => (x"7f",x"7f",x"7f",x"7f"),
    22 => (x"1c",x"08",x"08",x"00"),
    23 => (x"7f",x"3e",x"3e",x"1c"),
    24 => (x"3e",x"7f",x"7f",x"7f"),
    25 => (x"08",x"1c",x"1c",x"3e"),
    26 => (x"18",x"10",x"00",x"08"),
    27 => (x"10",x"18",x"7c",x"7c"),
    28 => (x"30",x"10",x"00",x"00"),
    29 => (x"10",x"30",x"7c",x"7c"),
    30 => (x"60",x"30",x"10",x"00"),
    31 => (x"06",x"1e",x"78",x"60"),
    32 => (x"3c",x"66",x"42",x"00"),
    33 => (x"42",x"66",x"3c",x"18"),
    34 => (x"6a",x"38",x"78",x"00"),
    35 => (x"38",x"6c",x"c6",x"c2"),
    36 => (x"00",x"00",x"60",x"00"),
    37 => (x"60",x"00",x"00",x"60"),
    38 => (x"5b",x"5e",x"0e",x"00"),
    39 => (x"1e",x"0e",x"5d",x"5c"),
    40 => (x"ec",x"c2",x"4c",x"71"),
    41 => (x"c0",x"4d",x"bf",x"d5"),
    42 => (x"74",x"1e",x"c0",x"4b"),
    43 => (x"87",x"c7",x"02",x"ab"),
    44 => (x"c0",x"48",x"a6",x"c4"),
    45 => (x"c4",x"87",x"c5",x"78"),
    46 => (x"78",x"c1",x"48",x"a6"),
    47 => (x"73",x"1e",x"66",x"c4"),
    48 => (x"87",x"df",x"ee",x"49"),
    49 => (x"e0",x"c0",x"86",x"c8"),
    50 => (x"87",x"ee",x"ef",x"49"),
    51 => (x"6a",x"4a",x"a5",x"c4"),
    52 => (x"87",x"f0",x"f0",x"49"),
    53 => (x"cb",x"87",x"c6",x"f1"),
    54 => (x"c8",x"83",x"c1",x"85"),
    55 => (x"ff",x"04",x"ab",x"b7"),
    56 => (x"26",x"26",x"87",x"c7"),
    57 => (x"26",x"4c",x"26",x"4d"),
    58 => (x"1e",x"4f",x"26",x"4b"),
    59 => (x"ec",x"c2",x"4a",x"71"),
    60 => (x"ec",x"c2",x"5a",x"d9"),
    61 => (x"78",x"c7",x"48",x"d9"),
    62 => (x"87",x"dd",x"fe",x"49"),
    63 => (x"73",x"1e",x"4f",x"26"),
    64 => (x"c0",x"4a",x"71",x"1e"),
    65 => (x"d3",x"03",x"aa",x"b7"),
    66 => (x"f7",x"d2",x"c2",x"87"),
    67 => (x"87",x"c4",x"05",x"bf"),
    68 => (x"87",x"c2",x"4b",x"c1"),
    69 => (x"d2",x"c2",x"4b",x"c0"),
    70 => (x"87",x"c4",x"5b",x"fb"),
    71 => (x"5a",x"fb",x"d2",x"c2"),
    72 => (x"bf",x"f7",x"d2",x"c2"),
    73 => (x"c1",x"9a",x"c1",x"4a"),
    74 => (x"ec",x"49",x"a2",x"c0"),
    75 => (x"48",x"fc",x"87",x"e8"),
    76 => (x"bf",x"f7",x"d2",x"c2"),
    77 => (x"87",x"ef",x"fe",x"78"),
    78 => (x"c4",x"4a",x"71",x"1e"),
    79 => (x"49",x"72",x"1e",x"66"),
    80 => (x"26",x"87",x"f9",x"ea"),
    81 => (x"71",x"1e",x"4f",x"26"),
    82 => (x"48",x"d4",x"ff",x"4a"),
    83 => (x"ff",x"78",x"ff",x"c3"),
    84 => (x"e1",x"c0",x"48",x"d0"),
    85 => (x"48",x"d4",x"ff",x"78"),
    86 => (x"49",x"72",x"78",x"c1"),
    87 => (x"78",x"71",x"31",x"c4"),
    88 => (x"c0",x"48",x"d0",x"ff"),
    89 => (x"4f",x"26",x"78",x"e0"),
    90 => (x"5c",x"5b",x"5e",x"0e"),
    91 => (x"86",x"f4",x"0e",x"5d"),
    92 => (x"c0",x"48",x"a6",x"c4"),
    93 => (x"bf",x"ec",x"4b",x"78"),
    94 => (x"d5",x"ec",x"c2",x"7e"),
    95 => (x"bf",x"e8",x"4d",x"bf"),
    96 => (x"f7",x"d2",x"c2",x"4c"),
    97 => (x"fe",x"e2",x"49",x"bf"),
    98 => (x"49",x"ee",x"cb",x"87"),
    99 => (x"cc",x"87",x"f0",x"cc"),
   100 => (x"49",x"c7",x"58",x"a6"),
   101 => (x"70",x"87",x"f3",x"e6"),
   102 => (x"87",x"c8",x"05",x"98"),
   103 => (x"99",x"c1",x"49",x"6e"),
   104 => (x"87",x"c3",x"c1",x"02"),
   105 => (x"bf",x"ec",x"4b",x"c1"),
   106 => (x"f7",x"d2",x"c2",x"7e"),
   107 => (x"d6",x"e2",x"49",x"bf"),
   108 => (x"49",x"66",x"c8",x"87"),
   109 => (x"70",x"87",x"d4",x"cc"),
   110 => (x"87",x"d8",x"02",x"98"),
   111 => (x"bf",x"ef",x"d2",x"c2"),
   112 => (x"c2",x"b9",x"c1",x"49"),
   113 => (x"71",x"59",x"f3",x"d2"),
   114 => (x"cb",x"87",x"fb",x"fd"),
   115 => (x"ee",x"cb",x"49",x"ee"),
   116 => (x"58",x"a6",x"cc",x"87"),
   117 => (x"f1",x"e5",x"49",x"c7"),
   118 => (x"05",x"98",x"70",x"87"),
   119 => (x"6e",x"87",x"c5",x"ff"),
   120 => (x"05",x"99",x"c1",x"49"),
   121 => (x"73",x"87",x"fd",x"fe"),
   122 => (x"87",x"d0",x"02",x"9b"),
   123 => (x"cd",x"fc",x"49",x"ff"),
   124 => (x"49",x"da",x"c1",x"87"),
   125 => (x"c4",x"87",x"d3",x"e5"),
   126 => (x"78",x"c1",x"48",x"a6"),
   127 => (x"bf",x"f7",x"d2",x"c2"),
   128 => (x"87",x"e9",x"c0",x"05"),
   129 => (x"e5",x"49",x"fd",x"c3"),
   130 => (x"fa",x"c3",x"87",x"c0"),
   131 => (x"87",x"fa",x"e4",x"49"),
   132 => (x"ff",x"c3",x"49",x"74"),
   133 => (x"c0",x"1e",x"71",x"99"),
   134 => (x"87",x"dc",x"fc",x"49"),
   135 => (x"b7",x"c8",x"49",x"74"),
   136 => (x"c1",x"1e",x"71",x"29"),
   137 => (x"87",x"d0",x"fc",x"49"),
   138 => (x"ec",x"c8",x"86",x"c8"),
   139 => (x"c3",x"49",x"74",x"87"),
   140 => (x"b7",x"c8",x"99",x"ff"),
   141 => (x"74",x"b4",x"71",x"2c"),
   142 => (x"87",x"dd",x"02",x"9c"),
   143 => (x"bf",x"f3",x"d2",x"c2"),
   144 => (x"87",x"c7",x"ca",x"49"),
   145 => (x"c4",x"05",x"98",x"70"),
   146 => (x"d2",x"4c",x"c0",x"87"),
   147 => (x"49",x"e0",x"c2",x"87"),
   148 => (x"c2",x"87",x"ec",x"c9"),
   149 => (x"c6",x"58",x"f7",x"d2"),
   150 => (x"f3",x"d2",x"c2",x"87"),
   151 => (x"74",x"78",x"c0",x"48"),
   152 => (x"05",x"99",x"c2",x"49"),
   153 => (x"eb",x"c3",x"87",x"cd"),
   154 => (x"87",x"de",x"e3",x"49"),
   155 => (x"99",x"c2",x"49",x"70"),
   156 => (x"c1",x"87",x"cf",x"02"),
   157 => (x"6e",x"7e",x"a5",x"d8"),
   158 => (x"c5",x"c0",x"02",x"bf"),
   159 => (x"49",x"fb",x"4b",x"87"),
   160 => (x"49",x"74",x"0f",x"73"),
   161 => (x"cd",x"05",x"99",x"c1"),
   162 => (x"49",x"f4",x"c3",x"87"),
   163 => (x"70",x"87",x"fb",x"e2"),
   164 => (x"02",x"99",x"c2",x"49"),
   165 => (x"d8",x"c1",x"87",x"cf"),
   166 => (x"bf",x"6e",x"7e",x"a5"),
   167 => (x"87",x"c5",x"c0",x"02"),
   168 => (x"73",x"49",x"fa",x"4b"),
   169 => (x"c8",x"49",x"74",x"0f"),
   170 => (x"87",x"ce",x"05",x"99"),
   171 => (x"e2",x"49",x"f5",x"c3"),
   172 => (x"49",x"70",x"87",x"d8"),
   173 => (x"c0",x"02",x"99",x"c2"),
   174 => (x"ec",x"c2",x"87",x"e5"),
   175 => (x"c0",x"02",x"bf",x"d9"),
   176 => (x"c1",x"48",x"87",x"ca"),
   177 => (x"dd",x"ec",x"c2",x"88"),
   178 => (x"87",x"ce",x"c0",x"58"),
   179 => (x"4a",x"a5",x"d8",x"c1"),
   180 => (x"c5",x"c0",x"02",x"6a"),
   181 => (x"49",x"ff",x"4b",x"87"),
   182 => (x"a6",x"c4",x"0f",x"73"),
   183 => (x"74",x"78",x"c1",x"48"),
   184 => (x"05",x"99",x"c4",x"49"),
   185 => (x"c3",x"87",x"ce",x"c0"),
   186 => (x"dd",x"e1",x"49",x"f2"),
   187 => (x"c2",x"49",x"70",x"87"),
   188 => (x"ec",x"c0",x"02",x"99"),
   189 => (x"d9",x"ec",x"c2",x"87"),
   190 => (x"c7",x"48",x"7e",x"bf"),
   191 => (x"c0",x"03",x"a8",x"b7"),
   192 => (x"48",x"6e",x"87",x"cb"),
   193 => (x"ec",x"c2",x"80",x"c1"),
   194 => (x"cf",x"c0",x"58",x"dd"),
   195 => (x"a5",x"d8",x"c1",x"87"),
   196 => (x"02",x"bf",x"6e",x"7e"),
   197 => (x"4b",x"87",x"c5",x"c0"),
   198 => (x"0f",x"73",x"49",x"fe"),
   199 => (x"c1",x"48",x"a6",x"c4"),
   200 => (x"49",x"fd",x"c3",x"78"),
   201 => (x"70",x"87",x"e3",x"e0"),
   202 => (x"02",x"99",x"c2",x"49"),
   203 => (x"c2",x"87",x"e5",x"c0"),
   204 => (x"02",x"bf",x"d9",x"ec"),
   205 => (x"c2",x"87",x"c9",x"c0"),
   206 => (x"c0",x"48",x"d9",x"ec"),
   207 => (x"87",x"cf",x"c0",x"78"),
   208 => (x"7e",x"a5",x"d8",x"c1"),
   209 => (x"c0",x"02",x"bf",x"6e"),
   210 => (x"fd",x"4b",x"87",x"c5"),
   211 => (x"c4",x"0f",x"73",x"49"),
   212 => (x"78",x"c1",x"48",x"a6"),
   213 => (x"ff",x"49",x"fa",x"c3"),
   214 => (x"70",x"87",x"ef",x"df"),
   215 => (x"02",x"99",x"c2",x"49"),
   216 => (x"c2",x"87",x"e9",x"c0"),
   217 => (x"48",x"bf",x"d9",x"ec"),
   218 => (x"03",x"a8",x"b7",x"c7"),
   219 => (x"c2",x"87",x"c9",x"c0"),
   220 => (x"c7",x"48",x"d9",x"ec"),
   221 => (x"87",x"cf",x"c0",x"78"),
   222 => (x"7e",x"a5",x"d8",x"c1"),
   223 => (x"c0",x"02",x"bf",x"6e"),
   224 => (x"fc",x"4b",x"87",x"c5"),
   225 => (x"c4",x"0f",x"73",x"49"),
   226 => (x"78",x"c1",x"48",x"a6"),
   227 => (x"ec",x"c2",x"4b",x"c0"),
   228 => (x"50",x"c0",x"48",x"d4"),
   229 => (x"c4",x"49",x"ee",x"cb"),
   230 => (x"a6",x"cc",x"87",x"e5"),
   231 => (x"d4",x"ec",x"c2",x"58"),
   232 => (x"c1",x"05",x"bf",x"97"),
   233 => (x"49",x"74",x"87",x"de"),
   234 => (x"05",x"99",x"f0",x"c3"),
   235 => (x"c1",x"87",x"cd",x"c0"),
   236 => (x"de",x"ff",x"49",x"da"),
   237 => (x"98",x"70",x"87",x"d4"),
   238 => (x"87",x"c8",x"c1",x"02"),
   239 => (x"bf",x"e8",x"4b",x"c1"),
   240 => (x"ff",x"c3",x"49",x"4c"),
   241 => (x"2c",x"b7",x"c8",x"99"),
   242 => (x"d2",x"c2",x"b4",x"71"),
   243 => (x"ff",x"49",x"bf",x"f7"),
   244 => (x"c8",x"87",x"f4",x"d9"),
   245 => (x"f2",x"c3",x"49",x"66"),
   246 => (x"02",x"98",x"70",x"87"),
   247 => (x"c2",x"87",x"c6",x"c0"),
   248 => (x"c1",x"48",x"d4",x"ec"),
   249 => (x"d4",x"ec",x"c2",x"50"),
   250 => (x"c0",x"05",x"bf",x"97"),
   251 => (x"49",x"74",x"87",x"d6"),
   252 => (x"05",x"99",x"f0",x"c3"),
   253 => (x"c1",x"87",x"c5",x"ff"),
   254 => (x"dd",x"ff",x"49",x"da"),
   255 => (x"98",x"70",x"87",x"cc"),
   256 => (x"87",x"f8",x"fe",x"05"),
   257 => (x"c0",x"02",x"9b",x"73"),
   258 => (x"a6",x"c8",x"87",x"dc"),
   259 => (x"d9",x"ec",x"c2",x"48"),
   260 => (x"66",x"c8",x"78",x"bf"),
   261 => (x"75",x"91",x"cb",x"49"),
   262 => (x"bf",x"6e",x"7e",x"a1"),
   263 => (x"87",x"c6",x"c0",x"02"),
   264 => (x"49",x"66",x"c8",x"4b"),
   265 => (x"66",x"c4",x"0f",x"73"),
   266 => (x"87",x"c8",x"c0",x"02"),
   267 => (x"bf",x"d9",x"ec",x"c2"),
   268 => (x"87",x"e5",x"f1",x"49"),
   269 => (x"bf",x"fb",x"d2",x"c2"),
   270 => (x"87",x"dd",x"c0",x"02"),
   271 => (x"87",x"cb",x"c2",x"49"),
   272 => (x"c0",x"02",x"98",x"70"),
   273 => (x"ec",x"c2",x"87",x"d3"),
   274 => (x"f1",x"49",x"bf",x"d9"),
   275 => (x"49",x"c0",x"87",x"cb"),
   276 => (x"c2",x"87",x"eb",x"f2"),
   277 => (x"c0",x"48",x"fb",x"d2"),
   278 => (x"f2",x"8e",x"f4",x"78"),
   279 => (x"5e",x"0e",x"87",x"c5"),
   280 => (x"0e",x"5d",x"5c",x"5b"),
   281 => (x"c2",x"4c",x"71",x"1e"),
   282 => (x"49",x"bf",x"d5",x"ec"),
   283 => (x"4d",x"a1",x"cd",x"c1"),
   284 => (x"69",x"81",x"d1",x"c1"),
   285 => (x"02",x"9c",x"74",x"7e"),
   286 => (x"a5",x"c4",x"87",x"cf"),
   287 => (x"c2",x"7b",x"74",x"4b"),
   288 => (x"49",x"bf",x"d5",x"ec"),
   289 => (x"6e",x"87",x"e4",x"f1"),
   290 => (x"05",x"9c",x"74",x"7b"),
   291 => (x"4b",x"c0",x"87",x"c4"),
   292 => (x"4b",x"c1",x"87",x"c2"),
   293 => (x"e5",x"f1",x"49",x"73"),
   294 => (x"02",x"66",x"d4",x"87"),
   295 => (x"de",x"49",x"87",x"c7"),
   296 => (x"c2",x"4a",x"70",x"87"),
   297 => (x"c2",x"4a",x"c0",x"87"),
   298 => (x"26",x"5a",x"ff",x"d2"),
   299 => (x"00",x"87",x"f4",x"f0"),
   300 => (x"00",x"00",x"00",x"00"),
   301 => (x"00",x"00",x"00",x"00"),
   302 => (x"00",x"00",x"00",x"00"),
   303 => (x"1e",x"00",x"00",x"00"),
   304 => (x"c8",x"ff",x"4a",x"71"),
   305 => (x"a1",x"72",x"49",x"bf"),
   306 => (x"1e",x"4f",x"26",x"48"),
   307 => (x"89",x"bf",x"c8",x"ff"),
   308 => (x"c0",x"c0",x"c0",x"fe"),
   309 => (x"01",x"a9",x"c0",x"c0"),
   310 => (x"4a",x"c0",x"87",x"c4"),
   311 => (x"4a",x"c1",x"87",x"c2"),
   312 => (x"4f",x"26",x"48",x"72"),
   313 => (x"5c",x"5b",x"5e",x"0e"),
   314 => (x"4b",x"71",x"0e",x"5d"),
   315 => (x"d0",x"4c",x"d4",x"ff"),
   316 => (x"78",x"c0",x"48",x"66"),
   317 => (x"db",x"ff",x"49",x"d6"),
   318 => (x"ff",x"c3",x"87",x"c8"),
   319 => (x"c3",x"49",x"6c",x"7c"),
   320 => (x"4d",x"71",x"99",x"ff"),
   321 => (x"99",x"f0",x"c3",x"49"),
   322 => (x"05",x"a9",x"e0",x"c1"),
   323 => (x"ff",x"c3",x"87",x"cb"),
   324 => (x"c3",x"48",x"6c",x"7c"),
   325 => (x"08",x"66",x"d0",x"98"),
   326 => (x"7c",x"ff",x"c3",x"78"),
   327 => (x"c8",x"49",x"4a",x"6c"),
   328 => (x"7c",x"ff",x"c3",x"31"),
   329 => (x"b2",x"71",x"4a",x"6c"),
   330 => (x"31",x"c8",x"49",x"72"),
   331 => (x"6c",x"7c",x"ff",x"c3"),
   332 => (x"72",x"b2",x"71",x"4a"),
   333 => (x"c3",x"31",x"c8",x"49"),
   334 => (x"4a",x"6c",x"7c",x"ff"),
   335 => (x"d0",x"ff",x"b2",x"71"),
   336 => (x"78",x"e0",x"c0",x"48"),
   337 => (x"c2",x"02",x"9b",x"73"),
   338 => (x"75",x"7b",x"72",x"87"),
   339 => (x"26",x"4d",x"26",x"48"),
   340 => (x"26",x"4b",x"26",x"4c"),
   341 => (x"4f",x"26",x"1e",x"4f"),
   342 => (x"5c",x"5b",x"5e",x"0e"),
   343 => (x"76",x"86",x"f8",x"0e"),
   344 => (x"49",x"a6",x"c8",x"1e"),
   345 => (x"c4",x"87",x"fd",x"fd"),
   346 => (x"6e",x"4b",x"70",x"86"),
   347 => (x"03",x"a8",x"c2",x"48"),
   348 => (x"73",x"87",x"f0",x"c2"),
   349 => (x"9a",x"f0",x"c3",x"4a"),
   350 => (x"02",x"aa",x"d0",x"c1"),
   351 => (x"e0",x"c1",x"87",x"c7"),
   352 => (x"de",x"c2",x"05",x"aa"),
   353 => (x"c8",x"49",x"73",x"87"),
   354 => (x"87",x"c3",x"02",x"99"),
   355 => (x"73",x"87",x"c6",x"ff"),
   356 => (x"c2",x"9c",x"c3",x"4c"),
   357 => (x"c2",x"c1",x"05",x"ac"),
   358 => (x"49",x"66",x"c4",x"87"),
   359 => (x"1e",x"71",x"31",x"c9"),
   360 => (x"d4",x"4a",x"66",x"c4"),
   361 => (x"dd",x"ec",x"c2",x"92"),
   362 => (x"fe",x"81",x"72",x"49"),
   363 => (x"d8",x"87",x"d4",x"d0"),
   364 => (x"cd",x"d8",x"ff",x"49"),
   365 => (x"1e",x"c0",x"c8",x"87"),
   366 => (x"49",x"c6",x"db",x"c2"),
   367 => (x"87",x"de",x"ec",x"fd"),
   368 => (x"c0",x"48",x"d0",x"ff"),
   369 => (x"db",x"c2",x"78",x"e0"),
   370 => (x"66",x"cc",x"1e",x"c6"),
   371 => (x"c2",x"92",x"d4",x"4a"),
   372 => (x"72",x"49",x"dd",x"ec"),
   373 => (x"dc",x"ce",x"fe",x"81"),
   374 => (x"c1",x"86",x"cc",x"87"),
   375 => (x"c2",x"c1",x"05",x"ac"),
   376 => (x"49",x"66",x"c4",x"87"),
   377 => (x"1e",x"71",x"31",x"c9"),
   378 => (x"d4",x"4a",x"66",x"c4"),
   379 => (x"dd",x"ec",x"c2",x"92"),
   380 => (x"fe",x"81",x"72",x"49"),
   381 => (x"c2",x"87",x"cc",x"cf"),
   382 => (x"c8",x"1e",x"c6",x"db"),
   383 => (x"92",x"d4",x"4a",x"66"),
   384 => (x"49",x"dd",x"ec",x"c2"),
   385 => (x"cc",x"fe",x"81",x"72"),
   386 => (x"49",x"d7",x"87",x"dd"),
   387 => (x"87",x"f2",x"d6",x"ff"),
   388 => (x"c2",x"1e",x"c0",x"c8"),
   389 => (x"fd",x"49",x"c6",x"db"),
   390 => (x"cc",x"87",x"dc",x"ea"),
   391 => (x"48",x"d0",x"ff",x"86"),
   392 => (x"f8",x"78",x"e0",x"c0"),
   393 => (x"87",x"e7",x"fc",x"8e"),
   394 => (x"5c",x"5b",x"5e",x"0e"),
   395 => (x"4a",x"71",x"0e",x"5d"),
   396 => (x"d0",x"4c",x"d4",x"ff"),
   397 => (x"b7",x"c3",x"4d",x"66"),
   398 => (x"87",x"c5",x"06",x"ad"),
   399 => (x"da",x"c1",x"48",x"c0"),
   400 => (x"75",x"1e",x"72",x"87"),
   401 => (x"c2",x"93",x"d4",x"4b"),
   402 => (x"73",x"83",x"dd",x"ec"),
   403 => (x"e4",x"c6",x"fe",x"49"),
   404 => (x"6b",x"83",x"c8",x"87"),
   405 => (x"48",x"d0",x"ff",x"4b"),
   406 => (x"dd",x"78",x"e1",x"c8"),
   407 => (x"c3",x"49",x"73",x"7c"),
   408 => (x"7c",x"71",x"99",x"ff"),
   409 => (x"b7",x"c8",x"49",x"73"),
   410 => (x"99",x"ff",x"c3",x"29"),
   411 => (x"49",x"73",x"7c",x"71"),
   412 => (x"c3",x"29",x"b7",x"d0"),
   413 => (x"7c",x"71",x"99",x"ff"),
   414 => (x"b7",x"d8",x"49",x"73"),
   415 => (x"c0",x"7c",x"71",x"29"),
   416 => (x"7c",x"7c",x"7c",x"7c"),
   417 => (x"7c",x"7c",x"7c",x"7c"),
   418 => (x"7c",x"7c",x"7c",x"7c"),
   419 => (x"75",x"78",x"e0",x"c0"),
   420 => (x"ff",x"49",x"dc",x"1e"),
   421 => (x"c8",x"87",x"d0",x"d5"),
   422 => (x"fa",x"48",x"73",x"86"),
   423 => (x"fa",x"48",x"87",x"ef"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

